-- Works in behavioral
-- Works in synthesized
-- FINE! (OK)

library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_11 is
end tb_11;

architecture project_tb_arch of tb_11 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
 
    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");
 
    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 32759;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      127,                                                        -- S
                                                      0, -1, 8, 0, -8, 1, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (51, 29, -5, -65, 1, 53, -17, -15, -3, -4, -17, -63, 73, 44, 17, 34, 35, 5, -2, 34, -35, -30, 13, -37, -56, 38, 41, -59, -18, -45, -28, -45, 59, 40, -35, -18, 17, 23, 40, -61, -59, -53, -51, -63, 67, 41, 46, 24, -31, -34, -17, 7, 11, 69, 45, 28, 29, 10, 44, -64, 38, -62, -34, 21, 53, 7, -74, -6, -48, 41, 6, -33, 64, 30, -21, 53, -6, -51, 1, 36, -10, 57, -33, 74, 49, -64, 24, 2, 19, -8, 13, -18, 3, 53, -75, -20, -18, -74, 47, 7, 43, -22, 49, 29, -70, -48, 6, -1, -24, -71, -41, 39, 62, -1, 35, 33, 10, -17, -41, -48, 48, 46, 7, -25, 23, 7, 28, -71, 7, 0, 11, -28, 53, -17, -75, 58, 10, 4, -20, 60, 6, 12, 21, -10, -64, -19, -53, 19, 37, -18, 46, 8, -48, -25, 58, 48, 58, 9, 52, -13, -67, -15, 34, 59, 41, 32, 39, -24, -42, -59, -42, 39, 29, 54, -46, 38, -43, -24, -19, 68, 33, -50, 0, 58, 0, -20, 30, -20, 64, 4, 42, 72, 63, -2, 53, 28, -46, 17, -74, -15, 33, -41, -51, -16, -64, -22, -54, -34, 27, 1, -42, -17, 26, 33, -35, -52, -64, 69, 4, 75, -3, -32, 70, -18, 42, 47, -67, 69, -14, -66, -21, -58, -33, 3, 1, -22, 54, 21, 17, 5, -54, 51, 63, 45, 6, -49, 66, 17, -56, -8, 15, 14, 36, 9, 70, 0, -20, -73, -9, 40, -64, 45, 57, -24, -30, -20, 29, -54, 74, -31, 25, -58, -56, 10, 62, 23, 36, 51, -35, 53, -33, 53, -8, -75, -14, -14, 0, 39, -14, 67, 3, -3, 34, -18, 49, -73, 38, 0, -52, 34, 44, 48, 52, 61, -17, 38, 9, -59, 13, 47, 70, 54, 22, -16, 54, -68, 43, -21, 46, -47, -32, -26, 23, 75, 29, -6, -74, -9, 70, -52, -50, 36, 69, 75, 20, -26, 37, -49, -9, -27, 71, -17, -49, 17, 42, -73, 24, 9, -19, -8, 35, 22, 39, -18, 22, -7, 52, 21, 57, 44, 44, -71, 2, 38, -72, -54, -64, 39, -28, 0, -64, -35, 58, -40, 57, 24, -38, 3, -45, 17, 71, 63, -37, 34, -30, 58, -51, -56, 4, -69, 63, -30, -65, -11, -70, -63, 9, -60, 51, 56, 15, 62, -56, -2, -56, -75, -56, -21, 2, -27, 71, -3, -40, -43, -47, 3, -63, -24, 22, 14, -18, 9, 60, -10, 72, 63, 2, 5, -73, -23, -17, 18, -39, 2, -62, -20, 1, -45, 33, -73, 1, 26, -3, 37, 56, 23, -36, 69, 74, 60, 5, -20, -7, -11, 44, -11, -25, -30, 67, -23, 23, -25, 68, 57, 52, -72, -40, -23, -41, 68, -23, 35, 18, 49, -6, -1, -5, 34, -10, -7, 18, 70, 47, -67, -18, 15, -4, 32, 60, -13, -67, 5, 35, 75, -13, 12, -73, 22, 62, -41, 12, -38, 70, -48, -65, -12, 26, 5, -56, -62, 72, 35, -67, 43, 42, -10, -18, -40, -56, -36, 20, -50, 43, -20, -51, -46, 67, -48, 49, 51, -14, -17, -63, -22, 10, -54, 40, -41, 24, 57, -28, 20, 15, -20, -15, -21, 43, 40, 14, 62, -71, -42, -63, 47, 13, -39, 74, 2, -14, 45, -24, 46, -48, -12, -54, 37, 7, 59, 71, -44, 41, -34, 49, -22, 21, -41, 32, -13, 74, -30, -27, -75, 1, -17, 47, -63, 18, 43, 14, -72, 12, 63, 47, 39, -24, 69, -1, 56, 52, -8, -64, 15, 33, 59, 68, -21, -58, 22, 41, -62, 65, -64, -61, -9, -5, 59, 3, -63, 27, -61, -62, -39, -73, 61, -75, -24, 52, -3, -44, 26, 64, -34, -36, 22, -51, -46, 74, -36, 52, 39, -25, 41, 48, -11, -44, -33, -29, 32, -23, 71, 45, -11, -46, 47, -26, -46, -55, -52, 24, -24, 47, 13, 15, -67, -41, 39, -37, -43, -73, -61, 69, -22, 55, 41, 40, -66, -69, -67, 41, -19, -74, 8, 45, -44, -21, -59, -17, -3, -38, -68, 47, -66, 20, -14, -58, 52, -50, -22, -67, -50, -8, -74, 1, -30, 40, -36, -21, 44, -28, -58, -50, -28, 26, 70, 3, -73, -66, 59, 0, -29, 66, -29, -22, 8, 32, -6, -16, 55, 47, -8, -70, -36, -9, 4, 9, -46, 43, 61, 73, -60, -73, -55, -13, 28, -62, 63, 31, -53, 46, -47, -7, 35, -3, 45, -33, -47, -37, 27, -69, -66, -59, -66, -29, 6, 13, 55, 35, -19, 40, 30, -6, 41, 49, 54, -9, 62, 41, -56, -69, 9, -28, -3, -32, 44, -34, 11, 71, 4, -40, -74, 12, -24, -65, 58, 55, 21, 36, 12, -74, -2, -35, -7, -37, -62, -29, 30, 73, -64, 49, -72, 21, -56, 0, 64, 63, 40, -3, 56, -32, 32, 57, 53, -69, 65, 36, 61, 11, -4, -2, 10, 69, 38, -72, -43, 51, -26, 60, 46, -16, 33, 49, -73, 52, -29, 64, 38, -67, -14, 18, -25, -58, -2, -48, -54, -15, 63, -68, 71, -17, 5, 4, -25, -35, 5, 7, -62, 54, -9, 59, -40, -54, 30, -38, 72, 74, -51, 32, -68, 10, -26, -18, 25, 45, 7, 47, -45, -5, 52, -52, 51, -19, 27, -50, 19, -46, 30, 32, -69, -57, 15, -34, -35, -33, 2, -41, -35, 26, 66, -30, -42, -38, 27, 56, -68, -43, 25, -40, 27, 1, -17, 0, 55, -67, 26, -2, -38, -22, -46, -32, -3, 42, 8, 37, -67, -68, 69, -26, 33, 57, 19, 64, -57, -31, 44, -52, 1, -8, -17, -50, 68, 40, 23, 48, 46, -29, -30, -70, 25, 0, -28, -54, -34, 55, 56, -27, 62, 49, 22, 17, 30, -37, 3, 46, 5, -31, 70, -70, 36, -25, -47, 29, -63, 52, 1, 58, -55, 44, 64, 45, -32, -42, 66, 8, -63, 44, 56, 72, 15, 0, 11, -33, 38, -62, -62, -32, -18, -70, -29, -57, -22, -2, 45, -9, -28, -30, -29, -8, -62, -43, -38, -20, -10, -50, 61, 0, 68, 39, -4, 7, -37, -71, 50, 74, -58, 61, -36, -2, 64, 9, 14, -34, -69, -17, 30, -24, 26, -74, 43, 37, -42, -73, -59, 24, -49, 75, -54, -57, 36, 18, 23, 72, 20, -5, 71, 36, -22, -43, -42, -34, 41, 47, 6, 45, -46, -40, -57, 55, -41, 62, 16, -9, 62, 31, -63, -65, 28, -42, -49, -11, 51, 50, -15, -6, -33, -22, -46, 21, 11, -13, 60, -26, -44, -10, -58, -17, 24, -40, -40, 56, -56, 49, -29, -69, 2, -17, -61, -45, 17, -34, 17, -10, -60, 75, 59, -20, -22, -63, -75, 62, -3, 61, -42, 28, -27, -27, -67, 70, 9, -32, 51, 28, -58, -54, 32, 17, 5, 45, 45, -56, -65, -14, 9, -52, -14, -9, 3, 37, 1, 4, 21, 74, -13, 52, 24, 33, -50, 31, 28, 34, 74, 3, -16, -62, 22, -61, 31, -51, 59, 0, -32, 67, 60, 51, -61, -32, -34, 17, -73, 42, -57, 23, 38, 3, -1, -15, -39, 24, -60, 64, -20, -62, -11, 38, -50, -65, 52, 56, -40, 33, -22, 1, 24, -38, -24, 36, 3, 17, -23, 5, -18, -6, -48, -56, 72, 25, 4, -45, -29, 19, -59, 27, 31, 5, -13, 56, 14, -39, 34, 47, 69, -66, -28, 15, -28, 24, -25, 50, -37, 25, -20, 20, -59, 5, 38, -64, -46, -34, -34, -1, 59, -19, -52, 14, 61, 10, -8, -3, 46, -50, -32, 37, -41, 14, -26, 4, -38, 22, -23, -2, -31, 30, -57, -14, -41, 56, -5, -13, -56, 36, 61, -73, -59, -67, 14, -75, 16, -70, -5, -14, -45, 37, -55, -12, -25, -6, 67, 10, -62, -32, -68, -18, 73, -52, 41, -45, -72, -40, 17, -52, 72, 0, -52, -65, 6, 38, -67, -54, 43, 4, 7, 72, -35, 25, -16, 13, -59, -27, -53, -46, 15, -46, 11, 10, -22, -23, 40, -21, 10, -21, 0, 6, 52, 24, 15, -18, -16, 21, 3, -49, -51, -68, -53, -13, 32, 4, 75, 48, 53, -54, 75, -10, -26, 11, 75, 25, 61, 38, -72, -5, -61, 2, 75, 67, -52, 12, -27, 7, -43, 52, 33, -20, 59, 54, 40, 14, -20, 40, -14, -45, 59, -16, 20, -45, 68, 18, 55, 51, -20, 57, -32, -6, -17, -35, -15, 6, 52, 34, -65, -68, 10, 43, -15, -9, 19, -51, -71, 75, 62, -11, -48, 46, 48, 48, -75, 40, -10, 54, 15, 43, 35, 58, -39, -60, -52, 20, 19, 73, -22, 29, -73, 61, -6, -13, -26, -62, 12, -21, -65, -2, 41, -40, -34, 13, -68, -33, -25, -5, -57, 63, -38, 53, 43, -3, 66, 64, -61, 9, 60, -8, -38, 62, -25, 29, -26, 24, 42, 59, -75, 50, -21, 41, -65, 21, -24, -60, 61, 24, 9, -72, 11, 46, 54, -23, -35, 44, -35, -21, -25, -51, 44, 10, -66, -59, -37, -17, 41, -72, -36, 39, 51, 18, 3, 61, -37, 54, 75, -54, 3, 8, -51, -64, -24, -75, -12, 17, 42, 29, 69, -59, 51, 36, 24, 58, 52, 63, -37, 15, 64, 2, -21, 39, -57, 57, 25, -19, 33, 24, 1, -40, -44, 25, -28, 5, 24, 33, -54, -10, -14, -62, 5, -40, 49, -47, -58, 25, -62, -19, -35, -74, 56, 17, 41, 74, -4, -12, -22, -47, -66, 54, -11, -37, 1, 34, 43, -51, -9, 63, 13, 51, -75, -58, -67, 49, -30, -52, -4, -16, 2, 34, -17, -17, -25, -52, -19, 44, 9, 34, 73, 18, 10, -16, 56, -64, -60, 24, -42, 6, 11, 46, -21, 11, 63, -15, -18, -44, 9, 53, 13, -65, 10, 71, -7, 60, -58, 48, 29, 26, 4, 24, -31, -61, -68, -51, -50, -53, 46, -19, 26, -19, -48, -72, 65, -63, -12, -29, -34, 72, -53, 54, -68, 32, 48, -2, 14, 63, -30, -35, 11, 48, 64, 55, 62, 69, -73, -66, -62, 46, -10, 38, -48, 15, 39, -61, 28, -49, -16, 69, -54, 6, 46, -49, -40, 16, 24, 47, 3, 68, -63, -64, 40, 74, 67, 24, 66, 67, 33, -74, 35, -55, 37, 60, 36, 0, 75, -14, 27, -17, -21, 46, 62, -53, 72, -56, 36, 18, 66, -39, 8, -75, -27, -30, 73, -38, 69, 61, -49, 26, 62, 61, 47, 24, 46, 7, -54, 45, 66, 46, -50, -31, 16, -64, -10, 12, -47, -52, -47, -57, -15, 36, -58, 33, -69, -61, 70, 75, 75, -57, 24, 59, -72, -7, 5, 49, 73, 27, 16, 63, -5, 39, -46, -64, 48, 17, 21, -75, 41, 47, -58, -50, 8, -41, 58, 12, -27, 50, 9, -30, 66, -43, -49, 69, 25, 30, 41, 20, -21, -21, 7, 49, -57, 37, 58, 66, -22, 4, 67, -57, -25, -67, -34, 56, -35, -54, -8, 11, 71, -74, 56, 59, -44, -71, 53, 55, 34, 18, -1, -63, 70, -71, 62, -63, 41, 44, -72, -59, -30, 68, -42, 19, -75, -1, -1, -35, 21, 65, 51, 14, 64, 29, -2, -56, 31, -27, 72, -10, 64, -4, 2, 58, 0, -14, 71, -37, -47, 72, -23, -2, 64, 8, -61, 62, -70, 14, -51, 26, 1, 73, -38, -11, 26, 33, 6, -21, -72, 3, 44, 67, 72, -31, 48, -6, 28, 43, 30, 56, 37, -71, -23, 25, 13, -9, 9, 18, -73, 33, -34, 1, 30, 1, 65, -22, -41, -6, 32, -40, 70, -1, -48, 66, 41, 75, -16, -7, 40, -64, -28, -1, -60, 24, -54, 28, -63, 30, -32, -62, -15, 9, 14, -61, -65, 2, -10, -33, 71, -56, 2, 65, 16, 27, 55, -19, 24, -39, 50, -14, -30, -54, 60, -15, 43, -70, -62, 53, 35, -21, 66, -58, 64, 5, -46, 72, -69, 19, -39, -74, 37, 38, 64, -23, -12, 41, 32, -64, 75, 4, -4, -31, 23, -20, 29, -10, -16, 40, -33, -59, -56, -44, -41, -70, 36, -12, -74, 42, -70, -38, 41, 42, 73, 27, -59, -17, -8, 48, -5, -9, -24, 64, 35, 74, -32, -12, -14, 27, -49, 27, 44, -30, 58, -75, -25, 18, -12, -26, -18, -7, 11, -55, -41, 6, 47, -26, 65, -39, -54, -18, 27, -4, -30, -16, -8, 13, 45, 52, -37, 71, 3, -71, -37, -15, -71, 11, -75, -8, 60, -20, 59, -5, -2, -58, 75, -33, -11, 64, 1, 9, -30, -50, -71, 13, 9, -6, -52, -24, -30, -14, -28, 48, -12, 8, -45, -10, -56, -47, 58, -72, 6, 39, -3, -72, 54, -4, -32, -32, -18, 44, 52, 25, 69, 56, -38, 0, -26, -15, 52, 18, 45, -54, -10, -45, 29, 21, 21, 48, 47, 1, 52, -22, -36, -29, -21, -58, 42, 23, -15, -54, -11, -41, 46, -17, -63, -70, 56, -15, -12, 32, -73, -45, 53, -8, -14, 7, -65, -69, -23, 58, 5, -49, -42, 44, -3, 12, 59, -39, -43, -33, -18, 22, 1, -50, -73, 14, -45, 58, 74, 17, 15, -75, 47, -10, -10, -43, 70, 1, -39, -28, -19, 39, -2, 14, 7, 69, -52, -9, -46, -19, 31, 10, -73, -44, 35, -73, 45, 64, 60, 41, 5, -3, 41, -24, 61, -44, 7, 55, 30, 41, -51, -65, 5, 21, 22, -66, 14, 45, -2, 43, -50, -47, -23, -50, -15, -65, -50, -48, 74, -65, 69, 3, 5, 32, 52, -10, 63, -19, -32, 17, -53, -8, 25, 25, -63, -31, 32, 26, -61, -45, -8, -38, -19, 42, -14, 39, 52, 11, 67, 48, 19, 60, -25, -51, 16, -50, 12, 2, 6, 55, -59, 26, -30, 40, -27, -18, -67, -70, -69, -55, -42, -4, -17, 14, -38, 42, -22, -63, -23, -31, 60, 70, -49, -42, -57, 40, -19, 28, -36, 60, 6, -19, 11, 51, -57, 57, -43, -49, 62, -39, -28, -58, 32, 28, 32, 68, -6, -68, -73, 44, -24, 62, 38, 0, -58, 54, -38, -2, 7, 2, -17, -63, 56, 67, 63, 74, 48, -58, -53, 33, -21, -6, 50, -67, -56, 4, 74, 13, 11, -75, -18, 60, 63, -58, -18, -73, 72, 20, 1, 3, -56, 57, 15, 73, 48, 0, 69, 18, 17, -60, -27, 69, 8, -54, -75, 27, 25, 74, -37, -41, 75, 18, -57, 60, 35, 1, 62, 31, -57, -15, -42, -40, -34, 46, -43, -64, -32, -50, 28, 59, -35, 74, 50, 46, -56, 50, -2, 45, 47, 36, -72, 46, -24, -56, 28, -65, 20, 14, 42, 36, 73, 73, 71, -39, 42, -48, -29, -68, -25, 74, 66, 16, 70, 41, -16, -61, 13, 57, 57, -16, 15, 58, -48, 66, -74, 55, 75, 20, -8, 39, -20, -11, 36, -26, 23, 0, 1, 69, 8, 50, 65, -4, -10, 60, -41, 47, 74, 48, 29, 55, -46, -34, 35, -20, -45, 36, -41, -46, -20, 24, 68, 34, -65, 26, -68, 34, -51, 6, 27, 30, -20, 17, -50, 43, 1, -15, 15, -3, -45, -34, -26, -16, 5, -67, 37, 35, 42, 72, 62, -55, 18, 52, 52, 29, 3, 57, -13, 25, -13, -62, -21, 41, 28, 4, 6, -47, 62, -57, 23, -59, -18, 70, -1, 63, -73, -40, 20, 43, -46, 5, 63, 48, -19, 39, 1, 57, 20, 63, 6, -71, 74, 60, 43, 27, -13, -28, 53, -27, -12, 1, -10, 46, -7, 62, 31, -6, -56, -25, -39, -26, 55, -54, -56, -41, 60, 20, -60, 2, 5, 22, 4, 3, 4, -30, -48, 66, 17, -70, -36, -71, 4, 27, 48, 72, 11, 3, -10, 30, 52, 26, -74, 29, 47, -55, 63, 29, 38, -72, -47, -35, 23, 31, 42, -49, -75, 69, -60, 15, 74, -23, 17, 2, -72, -10, -3, 12, 66, 62, -34, 42, 11, -34, -4, -20, -16, -17, -68, -53, -16, -40, -15, -71, 66, -49, -46, 64, -55, -31, 3, -59, 21, -55, 17, 22, 8, -62, -42, -2, 73, -3, -35, 8, 38, 36, 62, -53, -59, 69, -33, -1, -49, 27, 3, -60, 52, 30, -72, 70, 74, 5, -65, 17, 23, 25, -37, -45, 38, -6, 28, 34, 67, 68, -34, 29, 26, -50, 51, 41, -57, -60, -38, -30, 43, 40, -17, 19, -7, -16, 11, -9, 64, 21, -69, 11, -29, -31, 41, -69, 39, -6, 40, 28, -16, -71, -19, -65, -46, -45, 49, -29, -30, -65, 14, -65, 48, 72, 27, -35, -20, -38, 30, -33, 57, 36, 53, -50, -73, 17, -44, 39, -65, 70, -9, -8, 72, 46, 0, -50, -75, -27, -6, -30, -17, -68, -21, -46, -72, -70, -8, -18, -32, -54, 24, -51, 55, -1, -26, 58, -60, 3, 19, -52, -3, -65, 16, -9, 56, -60, 15, 54, -11, -67, -54, 45, -59, 0, 72, -58, 6, -11, -3, 49, 10, -55, 71, -10, 20, -31, -30, 35, 45, 64, 57, -35, 72, -3, 31, 52, 12, -30, 28, 74, -21, 50, 44, -7, -26, 40, 10, 53, -47, -68, 26, 37, -50, 19, -51, 43, 61, -6, 1, 31, -18, -18, 71, -23, 54, 24, -47, -10, 70, 55, -13, -29, 29, -45, 39, -75, 68, -29, 54, -56, -24, 2, 56, 2, -54, -71, -31, -69, -4, 43, 35, 51, -51, 28, -48, -73, -23, -21, -9, -31, -42, 53, 15, 60, -70, -24, 60, 73, 22, 38, -61, 74, -35, 68, -2, -14, 70, 40, -10, -10, 8, -50, -34, 30, 53, -9, 33, -48, 45, -54, -4, -75, 74, -65, 60, -74, -14, 45, 72, -69, 5, -64, -73, 45, -72, -2, -47, 74, -38, 19, -14, 43, 42, 27, -2, 17, -59, -47, 45, 61, -26, -35, 60, -30, -24, 44, -29, 35, 11, -33, 41, -59, -24, 41, 61, -20, -37, -63, -24, 1, 29, 37, -34, -5, -13, 39, -66, 3, 67, 54, -14, -37, -58, -30, 8, -9, -63, 52, -50, 23, -58, 65, 39, -7, 30, 23, 46, 69, 35, -54, -8, -12, 57, 31, 56, -32, -5, 65, 44, -16, 42, -46, 21, 59, -2, -49, -26, 10, -72, -1, -43, -55, -14, 70, 11, -61, 17, -18, -68, -24, 1, -3, 39, -18, -48, 17, 25, 20, 6, -9, -73, -28, 19, 23, -47, -59, 49, 2, 24, 50, 75, 54, 68, -15, 48, 4, -3, -11, 59, 4, 40, -16, 74, 1, 40, -51, -60, -13, 44, 22, 54, 46, 67, -3, -9, -55, 11, -37, 20, -41, -63, 19, -63, -70, -73, 61, 7, -1, -28, -10, -74, -65, 47, 73, 9, 11, -54, 25, 74, 66, -31, 52, 34, -40, -29, -52, -22, 57, -14, 74, -62, -4, 15, -52, -1, 15, -67, -70, -61, -21, -7, -62, -11, -37, -65, 73, 49, -43, 22, 45, -55, 66, 19, 52, -51, 65, 75, 2, 44, -17, -2, 57, 55, -64, -70, -22, 26, -64, -18, 40, -10, 50, 53, 52, -63, 62, 50, 60, -57, -6, 29, -39, -17, -27, -63, 7, -40, -65, -69, -71, -7, 3, 61, -30, 14, 64, 24, -36, 74, -70, -73, -12, 53, 53, -35, 64, 39, -63, 48, 57, 4, -1, -58, 62, 47, -47, -7, -68, -37, 0, -66, 29, -73, 68, 75, 14, 57, 23, 53, 55, 26, 55, -35, 1, 33, 3, -11, -4, 13, -41, -24, -58, 34, -9, -72, 3, 19, -3, 8, 55, 70, 17, 9, 70, 10, 8, 6, -11, -47, -17, -34, 52, -39, 4, -23, 69, -70, 40, -13, 18, 74, 36, 35, 30, -48, 37, -42, 44, -44, 41, 22, -52, -19, -47, -60, 64, 34, 21, -23, 60, -72, 16, 36, -36, -58, -65, -45, -53, 48, 16, 41, 47, -24, -2, 1, 1, -41, 32, -32, -12, -2, 63, 11, 54, -60, 26, 40, 49, -29, -59, 33, -27, 30, -9, 12, 47, -1, 41, 70, -28, -21, 33, -59, 30, -45, 15, -46, -12, -28, -5, 49, 43, -18, -15, 19, -5, -67, -17, -34, -20, -3, 72, 28, -49, -13, -38, 71, 59, -75, 63, -47, -21, 20, -31, -68, 49, 58, -41, -41, -48, 29, -68, 68, -67, -10, 11, 1, -1, 67, 42, 52, -12, 38, 4, 12, -53, 39, 5, -72, 38, -7, -43, -59, -63, -1, -52, 59, -19, -20, -58, 6, -67, -50, -2, -61, 15, -67, 15, -62, 73, -19, 65, -17, -59, -9, 68, -37, -47, -2, -33, 66, 64, -3, -71, 74, 71, -49, 58, -23, 6, 75, 56, 15, -51, -21, 27, 38, -15, -33, 49, -17, 21, 37, 39, 36, -48, 32, 74, -22, -48, -37, -34, -60, 33, -29, -62, 29, -3, 71, -72, -73, 71, 59, 15, -58, -38, -33, 53, 23, 7, 27, -72, -48, -12, 42, 63, 13, -4, 60, 67, 23, -55, -43, 38, 52, 1, 50, 5, 73, 43, 8, -75, 36, -11, 13, 54, 25, 55, 29, -30, -16, -20, -27, 10, 43, -63, -5, -21, 9, -23, -30, -44, -2, 0, 68, -26, 75, 42, 52, 72, 7, -18, 70, -32, 46, 8, -56, -5, -15, 48, 40, 45, -47, -65, -23, 69, -52, 47, -28, 32, -51, 15, 61, 20, -62, 53, 67, -63, 17, 43, -69, -53, -53, -74, -10, 66, 7, 9, -16, 65, -21, -54, 32, 5, -43, -67, -1, -22, 56, 44, -68, -73, -18, 68, 22, -7, 44, 11, 5, -17, -22, 9, 5, -2, 8, 68, -12, -61, -1, 47, -73, 54, 69, 34, -17, -50, 41, 55, 1, 19, 22, 8, 21, -74, 0, -35, -6, -34, 51, 72, 23, -49, 5, -48, 24, -62, -57, -64, -50, 17, 57, -48, -5, 50, 60, 52, 73, 23, 29, -2, -34, -27, -70, 60, -26, 3, -53, 41, 45, 71, 37, -8, -54, -35, 17, 43, -24, 35, 52, 1, -23, 33, 27, 45, 7, 9, 19, 2, -44, -29, 75, -5, 17, -73, -23, 65, 6, -1, 30, -27, -6, -10, 38, 13, 28, -21, -20, -72, -63, -46, 2, -13, 63, -49, -46, -8, 35, 49, 70, 64, -58, 67, -19, 34, 70, 31, 23, -2, -46, -24, 46, 21, 39, 8, -44, -9, 62, 11, -6, 72, 39, 69, -17, 26, -55, 13, -60, 53, -16, -68, 40, 1, 75, -57, -43, 67, 50, 54, -11, -72, -46, -43, 23, 66, 40, 54, -19, 24, -12, 48, 21, -49, 41, -74, 50, 59, 14, 63, 37, 73, 71, -1, -2, 68, 17, 29, 59, -9, 7, -30, -7, 34, 2, -60, 24, -36, 67, -71, 61, -23, 50, 4, 1, 15, 6, -27, -1, -56, -39, -42, -58, -44, 32, 13, -52, -27, -34, -71, 40, 46, -28, -43, 4, 49, -30, -50, -65, -41, -48, 71, 12, -74, 0, -65, 17, -70, -16, -62, -51, 20, -31, -36, 51, -75, 53, 72, -29, -59, 74, -67, 63, -30, -37, -11, -57, 8, 15, -49, 41, 42, -54, -25, 44, 19, -15, -17, 24, 44, -6, 47, -14, 38, -67, -39, 36, 59, -45, -69, -75, -47, -60, 61, -2, -24, -28, 14, 60, 62, 38, 23, 27, 60, 73, -5, 1, -20, 51, -50, -51, -33, 70, 10, -73, -75, 45, 38, 60, 73, 42, 58, -49, 55, 43, 22, -44, -61, -41, -62, 75, 72, 36, 26, 54, 31, -57, -20, -65, 67, 3, -43, -42, -5, 41, -40, -5, 8, 71, -21, 5, 37, -39, 29, 15, -74, -26, 46, -61, 6, 57, -64, 2, 17, 37, -21, -30, 53, 34, -20, 42, -41, 11, 75, 29, -24, -43, -52, 57, -48, 1, -14, 62, 35, -62, -1, 35, -13, -31, 49, 68, -52, 60, -8, 38, 19, 46, -68, -6, 2, -14, -40, 36, 72, -43, -11, -30, -11, 11, -49, 14, -64, 10, -2, 44, 21, 73, 3, -70, -36, -26, 71, -12, -44, -12, -50, 50, -44, -42, -34, 34, 17, 1, -6, 11, 31, 57, 56, -56, -8, -71, 31, 1, 12, -46, -31, -42, -49, 46, -37, -10, -56, -41, 53, -24, 20, -74, -52, 51, -41, -10, 7, 49, 64, -74, -16, 20, 58, -38, 37, -28, -34, -7, 48, 51, 22, -61, -69, 46, 60, -32, -42, -71, 0, -66, -22, -56, -65, 1, 68, -33, 64, 0, -60, 53, -1, -3, -5, -21, 34, -44, 26, 73, 24, -4, 48, -32, 10, 53, -64, -7, -55, -30, -5, 20, -23, 48, 39, -13, -29, 29, 27, -40, -47, 40, -65, 27, -39, 5, -70, 70, 36, 29, 67, -17, -51, 37, 24, 33, 14, 36, -50, 34, -72, 20, -24, -20, -10, -61, 40, 36, 44, -11, 69, 70, -47, -72, 22, -11, 6, 25, -19, -35, -21, -30, 23, 3, -69, -31, -40, 19, -73, -17, -25, -72, -75, 27, -19, -10, 39, -55, -51, 7, 7, -60, 0, 35, -56, -54, -54, 23, 44, 2, 63, -53, 47, 8, 26, 52, 53, 59, -7, 55, -35, 43, 57, -35, -6, -38, 29, -42, -19, 51, 38, 63, 66, -38, 21, -68, -19, 42, 31, -50, -31, 18, -30, -62, -49, 69, 63, -72, 53, -20, 56, -58, -52, 35, -20, 15, 73, -67, 46, -22, 59, 7, -37, 50, 42, 59, 57, -52, 26, 10, -29, 68, -47, 16, -72, -23, 10, 67, -20, -15, -29, -42, 0, -6, 69, 55, -68, 64, 62, 53, -36, 45, -16, 2, 17, -49, -16, -1, -28, -68, -69, 18, 73, -41, -44, -75, 11, 39, 67, 64, -54, -39, -55, 21, 30, -64, -1, 37, 75, -15, 13, -37, -46, 72, 38, 47, -53, -54, -32, -6, -47, -26, -66, -50, 7, -34, -51, -60, -71, -60, -71, -51, -26, -53, 45, -71, -42, -32, 39, -43, 26, -24, -7, 54, -29, -45, 25, -7, -25, 66, 61, 1, -38, 70, 27, 42, -40, 49, 58, -37, 62, 60, -13, -39, -69, -46, -37, -38, -4, -74, -6, -54, -24, 60, 75, 22, -61, 22, -63, -13, 10, 73, 64, 48, 68, 15, 14, -50, -14, -6, -14, -28, -22, 46, 8, -18, -75, 46, 19, -6, 46, -65, 15, -56, 70, 13, 41, -68, -43, 51, -6, 43, 47, -18, 13, 37, 70, -51, 62, -20, 19, -29, 28, 70, -59, -42, -23, -61, -71, 71, 8, 50, -71, -54, 69, 74, 32, 32, -70, 64, 5, -2, 29, -24, 53, -34, -63, 48, -11, 73, -50, -68, -32, 51, 75, -16, -66, -24, -1, -62, -30, -71, 61, -26, -50, 52, -30, 57, 6, -26, 46, -65, 45, -3, -15, 22, 39, -3, -6, -50, -8, 18, -45, 35, -7, -46, -58, 0, 4, 14, 11, 47, 18, -4, -57, 42, -30, -12, 23, 51, 35, -9, 60, 4, 64, -31, -49, 25, 39, 18, 50, -44, -40, -71, 64, 27, -44, -72, -49, 35, 17, 36, 6, -42, -46, 24, 75, 0, -65, 20, -27, 45, -64, -45, -28, 73, -1, -2, 22, -39, -62, -6, -10, -26, -2, -24, 74, 27, -20, -53, -13, 70, 58, 66, -50, -63, 13, -51, 10, 21, 43, 58, -12, 54, -62, 35, 51, 10, -45, -5, 44, -31, 64, -42, 16, -16, 10, 14, -65, 63, 34, -5, 55, 17, -16, -70, 29, 70, -48, -39, 15, 70, -57, -75, 46, -46, 34, 21, 40, 64, -62, 8, -43, -74, 40, 46, -17, -28, -18, -8, -43, -59, 62, -64, 31, -32, -59, -18, -38, -31, 18, 50, -37, 36, 51, -68, 66, 9, 26, 28, -5, 40, -42, 26, 39, 71, -4, -53, -33, 54, 14, -1, 68, -2, 9, 23, 42, 25, -71, -74, 67, 22, 50, -45, -20, 23, -40, -32, -44, 61, 71, 24, 25, -48, -26, -11, -53, 44, 9, -12, 20, -53, 62, 12, 20, -5, -43, -16, -57, -39, -14, -66, 56, -40, -38, -42, 56, -3, 2, -66, -17, -5, 33, -68, 22, -70, -6, 45, 49, -73, -43, -7, -53, -59, -73, 43, 10, -41, -51, 28, -7, 8, 35, -29, 41, 73, 4, 21, -8, -70, 30, 50, 1, -12, 56, -53, -7, -28, 65, -36, -25, -56, 32, -3, -39, 32, -38, 44, 64, -13, -6, -19, 68, -47, 27, 34, -52, -47, -21, 16, -41, -68, -12, 33, -5, -32, 53, 61, 16, 43, -51, 64, 62, 54, -17, -55, 10, 21, 62, -2, -70, -20, 52, 73, 7, 1, 29, 30, 29, -67, -32, 61, -60, 32, 18, 8, 73, -4, -9, 11, -39, 15, -1, -55, -9, 58, -36, 74, 1, -50, -6, 6, 6, -30, 1, -63, 44, -45, 40, -3, -39, -67, -19, -26, 38, 74, 55, 35, -8, -30, -29, 28, 58, 43, 47, -27, 23, -65, -31, -52, -40, 38, 27, 41, -70, -47, 51, 49, -19, 16, -32, 17, 22, 24, 66, -16, 21, 45, -59, -63, -63, -13, 39, 70, -47, 8, -35, 51, 18, 9, 73, 51, -31, 24, 15, -26, 50, -10, -55, -45, -72, -14, 47, 25, -67, 35, -69, 29, 2, -52, 39, 14, 8, 0, 6, 36, -70, 46, 10, 23, -21, 7, -1, 23, -47, -62, 70, -72, 1, -63, -44, 3, -1, -74, -50, 7, 36, -43, -42, -39, -22, 70, 48, 61, -7, -21, 20, -2, -51, -48, -56, 2, 32, 16, -53, 60, 27, -58, 61, -48, -46, -58, 30, 26, -57, 56, -45, 52, -65, -14, -65, -12, -21, 59, -29, 47, -40, 64, -33, -18, -60, -16, 59, 47, 75, -69, 30, 26, -54, 15, 52, -25, 30, 4, -74, 46, -18, -46, 23, -10, 16, 31, 53, 70, 12, -53, 41, 47, -65, -70, -46, -49, -10, -65, 71, -13, -59, 25, -64, -38, -37, 63, 11, 68, -11, 10, 39, 47, 39, -16, -39, -21, -61, -63, -29, 25, -41, -66, -4, -33, -60, 23, -9, 3, 34, -13, 63, 48, -64, 74, -67, -26, 59, 17, -33, -27, -49, -72, -58, 63, -13, -22, -35, -1, -12, 11, -52, 20, 21, 18, 63, 34, -37, -22, -39, 72, 38, -52, 43, 50, -55, 51, -54, -72, -10, -14, -24, 14, -11, -7, 1, 49, 45, 39, -29, -45, -25, -8, 51, 69, -68, 36, 27, -29, -64, 61, -35, 50, -67, -68, 22, -47, 56, 41, -45, -32, -48, 6, 57, 14, 75, -19, -14, 42, -56, 32, 72, -8, -54, 45, -15, -46, 3, -64, 0, 15, 72, 38, -13, -72, 44, -69, -46, 24, 47, -16, 68, 72, 64, 47, 11, 61, -48, 72, 27, -28, 26, 21, 39, 47, -9, -51, 74, 69, -42, -4, 6, -47, -41, 66, -46, -73, 70, -17, 24, 40, 41, 14, 36, 27, -16, -31, 12, 11, -35, -37, 58, 64, 57, 20, 34, -28, 42, 30, -36, 75, -49, 43, -48, -17, 32, -21, -17, 24, 36, -71, -12, 1, 17, -51, -48, -75, -7, 37, 11, 32, 73, -8, 18, 54, -64, -24, -51, 53, -69, -14, 50, -45, -49, -75, 13, 58, -21, 69, 7, -61, 73, 68, 13, 14, -59, 38, 12, 8, -1, -52, -36, -4, 13, 57, -25, 22, -44, -3, -3, -40, 58, -29, -10, -67, -31, -75, 65, 24, 69, -6, 36, 64, -14, -26, 1, 3, -66, -63, -65, 9, -42, -28, -73, 46, -49, -25, -8, -20, 47, 64, 15, 29, -42, -73, 36, 2, -73, 25, -52, 69, -57, 60, 56, 2, -44, -19, -71, -35, -9, -63, 47, 23, -18, 50, -7, 9, -51, 59, 62, 70, 45, 2, 21, -73, 4, -19, 5, 5, -72, 26, -4, -56, 10, -24, 22, 41, 30, 24, -71, -56, 37, 51, 42, -59, 23, -41, 23, 48, -60, 10, 40, 61, -64, -15, 63, 13, 40, -10, -60, 43, -59, 12, 61, 24, 61, 7, -12, 16, -45, -8, 35, 65, -35, -1, -69, 64, 33, 27, 36, 49, -39, 0, 32, -30, 58, 19, 57, 22, -68, 72, -10, -52, 8, -25, 47, -6, 55, -41, -68, -68, 24, 40, 73, 65, -37, -74, 53, 69, 26, 11, 40, 63, -67, -4, -45, 66, -62, -64, 13, -55, -67, -75, -32, 16, -27, -63, -68, -48, -28, -63, -41, 71, 52, -46, 60, -63, -47, 35, -69, 55, -30, 46, 40, -22, -35, 70, -31, -22, -69, 57, -2, -61, 55, 39, 28, -48, 51, 34, -21, -53, 46, 11, -59, 21, 41, 74, 33, 67, 34, 37, 46, -72, 6, 8, -20, 46, 3, 24, -54, 9, 3, 19, 23, -18, -18, -27, 9, -43, -69, 61, -22, 53, -4, -8, -4, -41, -10, -49, -51, -52, 62, 70, -50, -8, 3, 5, -40, -72, -49, -19, 12, 27, 73, -43, -67, -21, 5, 15, 9, 12, -2, 60, -13, 67, -24, 56, -49, 42, -69, -25, 63, 68, -33, -65, -18, 43, 15, 17, 46, 39, 71, -20, -10, 68, 12, -4, -31, -60, -65, 52, 25, 6, 36, -64, -2, -65, 65, 22, 50, 69, 70, 37, 60, -39, 48, -34, -73, -15, 57, 46, -51, 50, -49, 14, 43, 36, -67, -66, 51, -57, 59, 0, 23, 18, 9, -55, 28, -4, 42, 2, -10, 36, -39, -26, 70, -69, 13, 70, -8, -6, 41, 14, -31, 65, -50, -66, 23, -42, -59, -1, -25, -75, 72, 73, 18, 4, -58, -32, 75, 57, 45, -11, 15, -72, 36, 7, -65, -26, 2, 0, 41, -35, -62, -66, -48, -39, -59, 50, -5, -42, -29, 43, -44, -32, 40, 49, 47, 55, -59, 44, 34, 59, -42, -27, 62, 69, 55, 70, -33, -21, -6, -67, 19, 5, -60, 46, 42, -45, 21, -41, -14, 65, 75, 17, -43, 39, -12, -74, 16, 2, 46, -28, -17, -74, 20, -33, 70, -3, -38, -40, 52, 31, -34, -5, -41, -21, -36, -75, 9, 58, -43, 70, 47, -44, 9, -73, 68, 70, -72, 6, -4, 47, 53, 52, 48, -3, -56, 41, 69, -19, -75, 43, -66, -36, -39, -34, 18, 0, -34, -48, -20, -4, -56, -49, 25, 27, -49, 17, 21, -45, -53, -60, 75, 75, 67, 48, -6, -67, 11, -14, -13, 11, -49, -5, 48, -13, 36, -10, 62, -75, 15, -36, -4, 35, -9, -54, -16, 17, 36, -71, 45, 59, -58, 45, 56, -68, 15, -27, -60, -50, 32, 3, 34, 58, 73, 6, -30, 33, 69, -46, 33, 9, -6, -48, -34, 58, -27, 25, -3, -69, 27, -35, 65, 45, -68, 44, 52, 20, -61, 67, 45, 46, -6, 1, 26, -11, -71, 69, -53, 73, -54, 53, 6, 13, -71, 47, -7, -25, -4, 65, -18, -52, -48, -31, 68, -43, -65, 42, 52, -53, 33, 19, 66, -50, -56, 17, 12, -54, 8, 32, -56, 29, 10, 25, -34, 12, -5, 34, 61, 66, 22, -35, -64, 49, 9, -74, -71, 18, 43, 56, 40, -1, 0, 31, 22, 17, -30, -42, 39, 53, 66, 56, 5, -2, 3, 46, -66, 73, 5, 68, 62, -51, -43, 73, 71, 40, 73, 75, -18, 38, 56, -56, -41, -22, 48, 56, 68, -60, -63, 29, 69, -75, 9, -4, -2, -63, -34, 5, -66, 44, -4, 69, 68, 28, 67, 64, -8, 62, 61, 49, 24, 39, 67, 59, -59, 39, 37, -68, 55, 49, 36, 46, 47, -32, -34, -33, -20, 5, 46, -13, -26, -34, -19, -36, 69, -30, -48, -14, -44, -64, -43, 53, 50, -52, 36, 67, 61, -2, 74, 38, -31, 32, 8, -59, 75, 47, -17, -23, -24, -47, 38, 25, -8, -59, 65, -14, -14, -61, 45, 15, -50, -74, -8, -75, -52, -49, 65, -69, 22, 61, 44, 66, 15, -26, -71, 15, -55, -14, 65, -4, 12, 27, -54, -71, 43, -67, -12, -49, -55, -43, 41, -29, -44, -44, -31, -23, -18, -42, -17, -72, -59, -51, 67, 31, -2, 70, -32, 18, -22, -42, -63, 65, 58, -44, 67, 24, -36, -21, 50, -16, 9, 14, 28, 41, 43, 72, -58, -53, -48, -1, -50, -34, 21, -61, 73, -56, -69, -35, 35, -16, -4, 47, -28, -21, -73, -37, -73, -36, 16, 50, 24, -51, -14, -26, 63, -47, -29, -72, -25, -4, 2, -2, 38, -53, 11, 35, -36, 17, 73, 75, -74, -8, 44, -29, 46, 47, 9, 46, -65, -53, 18, 32, -28, -71, -69, -41, -45, -25, -38, 6, 46, 37, -74, 6, 58, 12, -37, -56, -46, -41, -57, -47, 26, 63, -1, -6, 32, -70, -36, 42, -47, 57, -3, -2, 59, 1, 30, -61, 51, 68, 18, 19, 27, 19, -50, 7, -44, -14, 27, -17, 20, 45, 11, -30, 30, -68, 39, -14, -65, -75, -49, -37, 56, 23, 36, 39, -54, -11, 51, 72, -19, -7, 13, -70, -63, 36, 13, -34, -53, -36, 24, 40, -69, -43, -65, 35, -38, 47, -55, -28, 48, -31, 9, 28, 65, -33, -11, -65, 31, -35, -71, -66, 31, 18, -60, 41, -24, 26, -69, -2, 63, 28, -37, 69, 58, -29, 28, -58, -58, 47, -10, 65, -60, 72, 15, -70, -37, -73, -62, 70, -35, -57, -72, 71, 34, -59, 35, -66, 42, 39, 6, 29, -8, 42, 21, -28, -63, -29, -10, -46, -58, 53, -58, -44, 49, 30, -41, -66, 32, -28, -74, 72, -12, -72, 66, -54, -56, 25, -46, 60, -12, 35, 11, 53, 1, -44, -50, 13, 3, 13, 40, 18, -12, 55, 49, -41, 8, -68, -32, -36, -22, -30, -41, 41, -27, -51, 61, -10, 47, -61, -28, -41, 47, 59, -63, -28, -63, -40, 58, 15, 46, 20, -44, -44, -2, -73, -10, -70, -67, 31, -33, -14, -75, 1, -51, -29, 23, -68, 35, -6, -56, -69, 27, 66, 65, 37, -40, -73, 72, -58, 15, 40, 36, 44, 71, -42, 47, -17, -37, 55, -62, 5, -37, -63, -71, -13, -19, 27, -5, -60, -54, 14, -55, 48, 3, -66, 9, 38, -66, 3, 56, 23, -35, 14, -11, -40, 47, -40, 16, -68, -61, 29, 10, -23, 41, 14, 38, -53, -36, -45, -38, -17, 44, -18, -47, -29, -10, 37, -68, -3, -38, 63, -58, 0, -1, 7, 33, -30, 42, -27, -25, 55, -74, 60, -46, 43, -3, 67, 63, 34, -54, -53, -59, 64, 3, -31, -43, 68, -72, -36, -13, -37, -51, 3, 38, 23, -66, -5, 66, 49, 43, -37, 26, 44, -54, 56, 9, 18, 45, -4, -24, 67, 17, -10, 53, -56, 34, -66, -66, 37, -28, -4, 75, -4, 72, 37, -58, -70, -46, -70, 53, 72, -31, 3, 38, -10, -17, -30, -70, -47, 41, -21, -58, -18, 44, 70, -1, 2, -74, 8, -39, -27, -73, -40, 43, 74, 70, 58, -73, -52, 63, 55, -58, -46, -18, 55, 19, 39, -51, 22, 67, 64, -75, -69, -32, 44, -75, 43, -32, 75, -27, 4, -29, -25, 37, -64, -26, 29, 69, -24, 50, 54, -45, 67, -69, 10, 45, 25, -27, 67, -28, -38, 55, -30, -32, -54, -63, -34, 62, -20, -34, -41, 58, 10, 10, 17, 21, 57, -31, 12, -45, -57, -10, -17, -67, -6, 68, 51, -56, -34, 42, -11, 1, 20, 32, 45, 41, 44, -67, 27, -53, -26, 59, -73, 59, -9, 19, 2, -28, 61, -62, 2, -73, 2, 60, -67, 71, 51, 59, -63, -61, 25, -1, 15, -31, -44, -16, -68, 75, -7, 32, -54, 40, 16, -52, 22, -71, 41, -54, -23, 26, -40, 52, 26, 35, 35, 34, 30, 10, 17, 41, 24, -35, -36, -37, 7, -5, 21, 15, -7, -64, -31, 12, 49, 60, 36, -7, 65, -1, 15, -36, -53, 48, -62, 49, 7, 48, 5, -41, -18, -53, 75, -72, -13, -38, -35, 67, 32, 61, 6, -53, 70, 51, 35, 41, 33, -7, -41, 20, 67, 49, 57, -64, 21, 71, 58, -50, 43, -12, -16, -52, 8, -16, -49, 68, 19, -11, 59, -25, -28, -12, -2, -34, -37, -45, -68, 69, 23, -34, 14, 12, -63, -7, 23, 31, -12, 4, 56, -46, 67, -36, -23, -3, 21, 1, -11, -36, 66, -28, 13, -38, 35, -67, 2, 71, -37, 9, 65, 61, 48, 1, -3, 58, 69, -58, 13, -20, 21, -7, 9, 10, 30, 59, -69, -24, -18, -5, 13, -30, 41, -50, 8, -2, -42, -68, -6, -4, 14, -19, -21, -16, 55, 49, -34, 46, 67, 54, -50, 10, -31, 32, -55, 74, 15, -51, -28, 73, 18, 61, -33, -17, -65, 48, 56, -33, 53, -28, 36, -9, 26, -60, 50, 5, 64, -62, -24, 53, 67, -1, -14, -42, -44, 4, -43, 44, 28, 4, 39, -30, -13, -71, 26, -2, 52, 7, 38, 30, 52, -2, -57, 3, 11, 67, -70, -2, -71, -19, -25, 72, 54, 34, -48, -68, -38, -16, 51, 66, 62, 15, -40, -27, 19, 62, 44, -7, -9, 6, -55, -35, -73, -38, 43, 13, -47, 47, -67, -43, -50, -16, -49, -72, -58, -21, -65, -20, 36, 60, -32, 22, -3, 3, 69, -62, -13, 35, 4, 51, -36, 25, -59, -34, 62, 57, 52, -63, 28, 61, -31, 54, -33, -6, 55, -18, 48, 64, 35, 8, 48, -73, -47, -31, 4, -54, -20, 64, 56, 59, 40, -58, 8, 54, -17, -8, 35, -42, 2, -14, -57, 47, -36, -17, -35, -59, 40, -65, -71, 0, 18, 52, 0, 44, -57, -72, 63, -2, 68, 42, -18, 32, 59, 63, 8, -35, -22, -33, -2, 55, 28, 14, 24, 65, 72, 64, -71, 34, 72, -67, -42, 13, 59, 32, -19, -74, 35, -31, -2, 27, -67, 55, -19, 67, 40, 64, -44, -58, -46, 27, 73, 55, -35, 21, 43, -41, 8, 47, 69, 4, 55, -51, -61, 38, 56, -4, 38, 14, 38, -40, -35, 46, -63, 20, 35, 52, 6, 67, 70, 35, 16, 65, 13, 57, 8, -20, -62, -62, -49, -71, 16, -72, -48, 30, 40, -68, -50, 2, 21, 61, 35, 60, 31, 47, 2, -9, 23, -70, -20, 15, 39, 71, 2, -24, 50, -67, 31, 62, -54, 55, 66, 37, 56, -58, -8, 20, -52, 15, -56, 42, 1, 54, 24, -46, 25, -50, 18, -29, -44, 73, 59, 70, 67, -14, -32, 39, -6, 72, 25, 13, 51, 14, -25, 29, 29, 40, -28, 52, -21, -9, 19, 55, -32, -33, -66, 68, -9, 25, -39, 22, 23, -55, 14, 12, 4, 57, -27, 71, 53, 72, 8, 26, 10, 56, -21, -37, 20, 24, -62, 75, -60, 32, 52, -17, 72, 59, -27, -13, 9, 8, -69, -46, 26, 18, 41, -46, -1, -64, -53, -26, -68, 28, 73, 15, 9, -23, 52, -49, 74, 65, -52, -62, 19, -75, -6, 13, 59, 41, -75, -10, -27, -71, 19, 74, 21, -18, -50, -56, -6, -28, -8, -1, 73, -11, -61, 4, 39, 66, 31, 38, 53, 54, 49, -4, 52, -32, -69, 36, -67, -71, -52, -21, -66, 43, -23, 30, -51, 2, 47, 16, 47, -39, -60, 42, 26, -46, -29, -11, -58, 75, -51, 68, 51, 74, -12, 28, -36, -8, -14, -28, -3, 9, 26, 6, -26, -75, -42, -1, 0, -73, -63, -29, -36, -48, -65, 65, -21, -19, -24, -4, -22, 1, -12, -48, -3, 49, 55, 36, -34, -37, -68, 38, 45, 31, -34, -56, 29, -3, 16, -47, -1, 28, -3, 36, 56, 7, 23, -43, 62, 73, 29, -36, -2, -61, -9, 70, 62, -32, 28, -50, 4, 33, 61, -26, -12, -51, -9, -61, 21, -69, -33, -58, 32, 39, 54, 10, -30, -1, 43, -46, -4, -6, -6, 67, 8, 58, 59, -8, -51, 11, 15, 26, -32, 0, 73, 29, 24, -12, 43, -33, -8, -66, -15, -53, 46, -39, 32, -61, 33, -1, -32, -46, 66, 35, -55, -3, 16, -71, 64, 38, 15, 4, -12, 59, -74, -14, 12, 26, 47, -22, 68, -38, -13, -25, -18, -44, 11, -62, -30, -31, 11, 13, -4, 1, -29, 16, 71, 62, 18, 60, 24, -44, -14, -66, -63, -13, -7, 24, -65, -37, 75, -72, -2, -13, -24, 55, 16, 63, 66, 61, -46, 1, -4, 23, -75, 42, -39, 71, 28, 55, 53, -26, -65, -39, -16, -53, 24, 50, 44, 34, -63, 44, 35, 10, -47, -64, -11, 44, 72, -20, 27, -52, 54, -53, 46, 52, 65, -69, 46, 15, 59, 23, 63, 69, 60, -31, -62, 6, -57, 58, -38, -44, 24, 73, 39, 50, -67, -47, 18, -73, 6, -33, -50, -18, -11, 69, -41, -24, 75, -71, 65, 59, 25, 52, 50, 7, -57, 64, -65, -39, 44, -27, -10, -10, -30, -46, -36, -24, -20, 55, -22, 59, -54, 1, -35, 8, -6, -1, 58, -9, 1, 47, -28, -51, 21, -53, 31, 39, -67, 42, 73, 52, -63, -12, -36, -18, 15, 3, 31, 68, -18, -69, 51, 1, 7, -60, -67, 74, 13, 66, -11, -62, 35, 37, -40, -20, 57, 65, -59, 65, 29, -61, 39, 41, 0, -73, -55, -63, 5, 51, -71, 60, 57, 55, -17, -14, 68, -9, -16, 5, -20, 46, 17, -61, 7, 52, -7, -12, 41, 9, -25, -6, 21, -62, -43, -57, -60, -23, -47, 18, -48, -43, 0, -69, -66, 58, -10, -73, -26, 49, 7, 27, 18, -52, 39, -51, 74, -44, 11, 37, 39, 59, -46, -18, 73, -14, 1, -65, 39, 27, 27, 64, 60, -49, 69, 67, -66, -17, 69, -19, -45, -1, -68, 48, 20, 46, 70, 16, -75, 3, -22, 39, -13, 7, -57, -18, 66, 17, -8, 27, -31, -57, 16, -49, -30, 7, -58, -23, 63, -66, 33, -58, 6, 38, 63, -50, 6, 58, 42, 4, -17, -58, -35, 43, 22, -16, -51, 12, -75, 17, -36, -31, 33, 53, -5, -75, -16, 11, -23, -29, 20, -68, -13, -50, 43, -26, -27, -26, -46, -63, 53, 13, -46, -57, -20, 51, 0, 3, -14, 0, -58, 25, 43, 50, 2, -40, 49, 59, 46, -52, -48, -12, -46, 14, 13, 72, 62, 60, -32, -60, 72, -54, 26, -51, -38, -71, 73, 37, 7, -17, -41, 24, -68, -74, -4, 7, -38, -31, -12, -70, -9, 16, -6, 20, -48, -69, 16, -62, 66, 60, -46, 61, -72, 53, -66, -37, 57, -69, 75, -14, -12, -44, -66, -5, -42, 6, -75, -7, 48, -12, -2, -37, -72, 67, 58, -44, 72, -3, -33, 60, -19, -6, 43, -16, -28, 52, 20, -49, 57, 17, 13, -31, 48, 22, 37, -72, -50, 35, -4, 72, -52, 68, -43, -51, 57, -60, -22, 51, 12, 21, 36, 66, -61, 3, -28, -16, -22, 67, 11, -43, 8, -54, -1, -20, 41, -42, -18, 65, 69, 51, 61, -59, 43, -58, -37, 23, -45, 17, -2, 40, -40, -44, 30, -28, 33, -74, 32, -65, 66, -35, -35, -2, -16, 39, 52, -51, 72, -42, -62, 65, -67, 72, -72, 50, -61, -33, -3, -33, 57, 70, -68, -59, -51, 37, -14, 57, 37, -58, 67, 27, -20, -46, -50, 37, 68, 75, 62, 62, -43, 73, 52, -35, 70, 53, -61, -69, -58, 9, -27, 74, 2, -22, -63, 26, -60, -1, 7, 50, 14, -4, 1, 68, 25, 24, 29, 15, 23, 13, 1, 55, 11, -23, -57, 5, -47, -45, 9, -30, 40, 55, -33, -34, -42, -23, 67, -27, 49, -4, -53, -14, 65, 21, -22, 14, -32, -71, -47, 66, 18, 29, 44, -49, -71, 62, 29, -45, -61, -38, -2, 54, -59, 38, -58, -26, -60, -69, 20, 62, 2, 40, -28, -9, -16, 23, -73, 27, 26, -47, 17, -34, 56, -17, -8, 58, -33, -55, -63, -18, -20, 10, -40, -4, -27, -22, 44, -14, -16, -14, -28, 60, -49, 18, -27, 10, -37, -24, -39, 64, 2, 51, -46, -18, -41, 19, -36, 1, 39, -24, 56, -59, 60, -59, 11, -45, -8, -21, 14, 49, 38, 61, 33, 64, 1, -71, -4, 40, -20, 30, 26, 55, 6, 54, -38, 38, -3, 1, -39, -41, 51, -58, -25, 33, -44, 61, 63, 23, -38, 1, -4, -75, -16, -48, 62, 61, -44, -17, 23, 9, -63, -29, -12, 16, -51, 25, -22, 22, -51, 13, 54, 73, 30, -47, 30, 61, -63, 17, 6, -28, -58, 75, -30, -1, -49, -43, -18, -20, 13, -71, 62, 25, -26, -27, -36, -2, 73, 15, -56, -56, -48, 71, -59, 55, -51, 46, 40, -41, -15, -32, 6, 0, -32, 50, 75, -8, -71, -19, 48, 17, -16, 32, -36, 33, -71, 3, -47, -75, -57, -29, -56, -32, -34, -41, -52, -10, -73, 63, 22, -12, -46, -49, 61, -3, -75, 60, 64, -71, -36, 34, 21, 21, -11, 58, -24, -7, -14, 4, -7, 2, 50, 11, 45, -61, 43, 68, 4, 45, 54, -51, -45, -68, -25, -59, 2, -25, 74, -12, -23, -40, -55, 71, 54, 9, 53, -46, -74, -39, 32, -7, 36, 4, -72, 6, 18, 44, -4, -55, 13, -28, -31, 44, -23, 17, 58, 54, 65, 56, -35, -34, -61, -15, -39, 68, 69, -64, -55, 68, -27, 52, -17, -67, -22, -16, 12, 70, -48, -69, -63, 41, -22, -21, 7, 31, 71, -11, 7, 60, -33, 47, -52, -19, -46, -16, -28, -55, -5, -8, -62, 41, -34, -6, 48, 17, 54, -18, 11, -70, -12, 23, 44, 40, 75, -27, -5, 70, 35, 75, 52, -73, 47, 75, -19, -75, -19, 26, -54, 50, -58, -43, 13, -17, 26, -15, -75, 2, 43, 9, 8, -47, -45, -26, 68, -46, 23, -15, -53, -18, -15, 72, -18, -46, 70, 37, -46, -25, -13, -27, -53, 3, 3, 36, 61, -48, -57, 59, 29, 59, -9, -41, -65, 21, 7, -73, 48, -46, -12, 68, 9, 46, 65, 65, 75, 57, 24, -49, -46, -65, 0, -23, 13, -75, -65, -3, -50, -49, -22, 55, -67, 42, -64, -57, -13, 18, -57, -42, 45, 6, -52, -21, -24, -65, -34, -25, 67, 65, 0, -54, 73, 75, -4, 11, 73, 4, -70, -52, 30, -19, -75, 36, -52, -64, 54, 8, 28, 71, 39, -3, 1, 63, 49, 51, 73, -61, -52, 65, -74, 23, -67, 75, 20, 4, 8, 16, -70, 11, 39, 33, 67, 39, -6, -61, 48, -30, 21, 0, -35, -16, 71, 40, -29, 44, 13, -31, 57, 36, -44, 58, -16, -38, 55, -74, 41, -13, 17, 44, 73, -22, 1, 65, -61, 70, -74, 63, -37, 20, -15, 3, -71, -20, -35, -25, -53, 53, 17, -74, 14, 46, 59, 71, -68, 39, 70, 46, -52, 12, 14, -54, 65, -60, -67, -73, -68, -68, 65, -30, 28, -28, 47, 32, 26, -64, -71, 46, 65, 20, 47, 1, -10, 28, -6, -2, -11, -12, -34, 13, 73, 56, 34, 61, 71, 40, 63, -73, 45, 50, -27, -3, -56, -58, -49, 45, -47, -44, 13, -60, 49, -16, 16, -37, -63, -68, 34, 1, -6, -75, -62, -9, 56, 45, -26, 49, 7, -39, 51, -23, -67, -54, 47, -47, -37, 74, 71, -10, -48, 9, 5, -75, 68, -56, -39, -73, -49, 71, 4, 20, 71, 15, -66, 49, -17, -17, 22, 63, 18, -5, -38, 26, 17, -66, 54, 53, -68, 50, -33, -43, -17, 48, -45, -27, 65, -9, -24, -60, -14, 53, 34, -21, -10, 41, -48, 46, -52, 49, 34, 41, -33, 71, -10, 59, -71, -32, 36, -66, -60, -74, -36, -4, 49, -6, 43, 38, 61, -57, 51, -29, 69, 7, 24, -17, -28, 51, -46, -6, 23, 61, -41, 65, 56, 22, 46, 59, 64, 4, 66, -72, 5, -45, -2, -24, 24, -35, -62, 7, -19, 63, 54, -26, -6, 2, 30, 40, -25, 57, -42, 73, 42, -10, 60, 23, -63, 30, 4, -75, -41, -6, -74, 39, 22, -1, -60, -31, 37, -49, 51, -58, -64, 27, -11, 6, -49, -58, -30, 2, 74, 1, -3, 41, 66, -18, -14, -73, -66, 65, -73, -34, -19, -71, -70, -72, 1, -57, -28, -39, -33, -53, -22, -21, 50, 41, 58, 74, 58, -50, 0, 56, 26, 71, 19, 16, -25, -71, 19, -16, 67, 21, 26, -27, 23, 29, -26, -53, 47, 21, -17, -64, 41, 34, -10, 13, -3, -28, 12, -21, -3, -66, -42, -53, -71, 50, 39, -21, 55, -18, 39, 44, -75, -13, -61, 22, -60, -12, 42, 60, -69, -51, 71, 46, 56, -14, -17, -22, 31, 68, 30, -47, -73, 63, -27, -71, 36, -66, -16, 13, -9, -55, -19, -10, 7, -4, -66, 20, 59, 51, 4, 64, 73, -3, 34, 53, 56, -61, -45, 10, -68, 61, 36, -68, 46, -67, -64, 6, -57, -7, -59, 7, 13, -2, 70, -58, 69, -72, 37, 50, 52, -37, 36, 47, 34, -6, 25, 14, 9, 53, -52, 16, 36, 59, 21, 7, 66, 32, -65, -67, -50, -48, 13, 36, 23, 8, 54, 14, 9, 15, -14, -16, 52, -53, -45, 10, 16, 53, -54, -51, 29, -32, 38, -11, -51, -17, 69, -61, -62, -73, -55, -39, -48, 34, 72, 50, -36, 50, -12, 48, -12, 49, -46, -36, 69, -17, 47, 10, -40, 68, 32, 64, -40, -5, -22, -15, 51, -31, -3, 64, -29, 18, -51, -2, -26, -56, -30, 13, 69, 33, -17, -19, 5, 13, 18, -2, 71, -11, -70, -47, -18, 38, -58, 15, -45, -7, 75, -70, 35, -3, 68, -69, -63, -61, 2, -14, -42, 48, 74, -50, 3, -21, 6, -70, 67, -51, 2, 60, 13, 7, -62, 68, -33, -47, 8, -3, 19, 5, 1, -22, 75, -7, -18, -64, 5, 60, -5, 39, 30, -9, 62, -45, 46, -8, -39, 35, 14, 38, 20, -50, -33, 31, -60, 10, 57, 23, -71, -2, -49, 5, 51, -50, 71, -44, -38, 1, -62, 32, -38, 43, -52, -52, 73, 67, 13, -44, 26, -48, 67, -32, -25, -41, 72, -10, 42, 51, -64, 44, -27, -38, -26, -53, -13, -31, -22, 22, 43, -9, -23, -71, -44, -2, -48, -49, -11, 39, -17, -63, 66, -26, -19, -37, 6, -25, 26, -28, -49, 37, -59, -1, 74, -12, 19, -16, 30, 72, -70, -2, -15, -20, 0, 16, 53, 28, 43, -34, -11, -52, -23, -21, -3, 33, 15, -72, -70, -35, -27, -44, -73, -13, 29, 74, 48, -28, -20, 3, -33, -14, -75, 27, 39, 0, -34, 17, -50, -69, 56, 14, -46, -43, 66, 26, 63, 3, 27, 69, 44, 74, -53, 44, -17, 49, 42, -44, -54, -53, 34, -12, 6, 32, -63, -31, -46, -22, 59, -22, -16, 40, 65, 13, 70, 54, -38, 58, -19, 62, 49, -51, 60, 69, 68, -34, 43, 33, -3, 62, 53, -47, -28, -19, 60, -16, 23, -64, 36, 7, -11, -56, -31, -21, 31, -39, -43, 66, -59, 11, 50, 65, 36, 33, 57, 26, 74, 24, -19, -5, 10, -42, 23, 55, 12, 5, -37, -42, 16, 72, 40, -72, -61, -69, -20, 45, -33, 10, 33, -16, -55, 7, -29, 56, -38, -48, 5, -40, 49, 61, 28, -19, -58, -27, -40, 27, 53, -3, 60, -8, -7, 22, -5, 7, 28, 48, -26, 69, -18, -71, -25, 2, 10, 19, -19, 47, 45, 59, -68, 18, 44, 33, 73, 59, -69, -43, 11, 59, 29, -5, -27, -53, -60, 41, 27, 41, 13, -74, 34, 70, -70, -69, -5, 15, 24, 49, -13, -7, 32, -8, -67, -2, -51, -70, -18, -45, -39, 66, -63, 65, -17, -15, -66, -2, -49, 37, -36, 39, 36, 71, 32, 39, -75, -51, -21, 24, 73, 39, -61, 29, -47, -53, -49, -23, -49, 6, 6, -13, -4, 18, -26, 55, -75, -18, -23, -51, -59, 14, 64, 52, 8, 18, 15, 8, 42, 67, -46, 39, 30, -32, -10, 58, -12, 16, -42, 12, -53, 37, 74, 16, -23, -27, -5, -23, 28, 46, 2, 44, -18, -12, 20, 65, -72, -43, -3, 45, -51, 26, 6, 52, 67, 69, 33, -22, 9, 66, 65, 29, 25, 64, -30, -74, -41, 38, -22, 62, 6, 53, 30, 64, -37, -28, 53, -34, 4, -27, -67, 28, 72, 12, 3, 64, 5, -40, -34, -63, -52, -45, 39, 48, -59, -67, 49, -27, 45, -51, -41, -25, -73, 62, -37, -37, -42, -61, 5, 36, -13, 13, -12, -19, -50, 64, -31, 28, -52, 8, 40, -29, 37, 4, -59, 51, 10, 65, -51, -21, -63, -17, 28, -63, -32, 64, -25, -1, -73, 55, -41, -13, -9, 21, 44, 14, 9, -65, -34, 33, 17, -69, -74, -24, 8, -57, -49, -60, -70, -25, -7, -58, 32, -55, -46, 75, -67, 5, -2, -66, -18, 33, -6, 48, -22, -40, -14, 62, -31, 28, 17, 61, 32, 19, -39, -38, 37, -13, -23, 42, 36, 45, 60, -8, 63, -64, -9, 72, 14, 64, -72, 72, 19, -5, 44, 70, 31, -47, 57, 75, 54, -4, 58, 8, -61, -59, 45, 49, 1, -56, 14, -39, 65, -2, 28, 52, 7, -59, 46, -54, -72, 47, -58, 22, -33, 59, 15, 71, -64, -4, 68, 65, 65, 48, -3, -71, 64, -36, 51, -13, -16, -11, 22, -29, 60, -26, -53, -8, -11, 67, 13, -8, 36, 28, -64, -75, 11, 26, 71, 21, -56, 61, 10, -66, 33, -70, -64, 19, -31, 62, -71, 28, -24, 26, 74, -40, 73, -56, 25, -14, -67, -38, 51, 42, 63, 61, 43, -3, 11, 36, -58, 29, 20, 27, 36, -23, 30, 47, 70, 75, 31, 74, 25, -69, 22, 22, -35, 19, 39, 65, -70, 45, -50, 54, 11, -63, 39, -22, 9, -25, -63, 26, -74, 32, -24, 37, -69, -70, 8, -75, -73, -37, 72, 28, -32, 18, -28, 8, -38, -65, -3, -35, 55, 22, -57, -10, 33, 58, 42, -36, -45, 54, 66, -46, 8, -36, 66, 14, -33, -4, 15, -32, 32, 9, 71, 75, -48, -35, 5, -13, -25, -75, 27, -48, 20, 43, 15, -23, 23, -21, 17, 51, -45, 5, -71, 38, 42, 70, -23, -67, -10, 65, -24, -55, -2, -31, -56, 23, 7, 23, -66, 55, 23, 34, -69, -33, 0, 20, 18, -53, 74, -43, 72, -46, 35, -75, 67, 1, 69, -34, 7, -19, -45, 57, 1, 29, -52, 21, -26, 31, -32, -16, 10, 64, -60, 15, -45, 15, -41, 46, 36, -43, -73, 32, -16, 37, 32, -26, -40, 23, 15, 43, -71, 44, 24, 5, -5, 47, -50, 44, 0, -9, -48, -65, -23, -34, 23, 6, 56, 57, -24, 14, -64, -23, -30, -6, -62, -75, 43, -26, 23, -20, -61, 27, -52, 36, -43, 18, 5, -20, -13, -70, 45, 12, -62, -54, 53, 36, 27, 32, 15, -74, -30, 26, -22, 14, -56, -11, 14, 60, 36, -41, -35, 50, 62, -14, 10, -59, -73, -62, -6, -11, -57, -39, 74, -46, -17, 50, 65, -68, 6, 4, -67, 49, -48, -14, -13, -30, 49, 74, -46, 9, -42, -8, -16, -58, 54, 67, -42, 56, -71, 25, -33, -55, 62, -37, -26, -33, -63, -39, -26, 16, 38, -17, -10, 66, 42, 50, -40, 15, 49, -13, -53, -71, 55, 6, -54, 31, -5, -23, 9, -2, 75, 49, 16, 61, -64, 66, -48, -53, -51, 0, 36, 63, 56, -50, 51, 22, 74, -67, -40, 45, -5, -18, 47, -28, 61, 68, -75, -22, -33, 9, 51, -34, -20, -8, -50, -8, -20, -23, 12, 4, 52, -28, -11, 32, -4, -36, -23, -6, -30, 10, -39, 41, 65, -68, -65, 48, 73, -64, -50, -36, 20, 75, 3, -75, -11, 28, -10, 44, -72, 75, -30, 53, -29, 33, 8, 42, 70, 58, -42, -35, -8, -8, -72, -21, -1, -62, -49, -6, -53, -26, 31, 41, -27, -41, 39, 37, 60, -47, 3, 61, -50, 47, 39, -4, 2, -31, -39, -4, -49, -8, 34, 16, 58, 37, 68, -21, 49, -57, 49, 69, -8, 4, 34, 39, 36, -3, -2, 21, 23, -74, 6, 48, 46, -33, -33, -28, 11, 3, 41, 35, 68, 0, -27, 50, -41, -35, -46, -70, -19, -73, 75, 49, 4, 33, 10, -35, -45, -68, 61, 51, -69, -11, 24, 50, 30, 66, -54, -37, -9, 61, 74, -19, -15, -31, -46, 17, 10, -17, 23, 64, -17, 22, 35, 62, -23, -31, -51, 7, -23, -68, -19, -19, -3, -71, -44, -49, 68, -25, -13, -19, -40, -17, 37, 18, 28, 66, -40, -40, -29, 56, -52, 29, 2, 59, 14, 54, -48, 38, -16, 2, 46, 40, 59, -35, 42, -63, -11, 34, -13, 51, -61, 23, -41, 49, -35, 60, 38, -2, -56, -67, -22, -33, 36, 53, -52, -26, 30, -26, -66, -62, 51, 53, 51, 32, -60, 15, 44, 4, -27, -44, -22, -15, 52, 10, -44, -61, -6, 69, 13, 13, -73, 66, 53, 36, 42, -74, -68, -4, -25, -59, 9, -52, 68, -18, 56, -70, 72, 22, 8, -33, 51, 61, 25, 27, -7, 54, 42, 62, 48, -23, -1, 48, -35, -26, 8, -69, -27, 15, 2, 23, 29, -67, 45, 19, -12, 23, 25, -18, -31, -43, 24, -57, -60, -29, 45, 8, -50, 9, -6, 71, 59, 66, 43, -53, -38, -27, -47, 11, 61, 29, -44, 14, 37, -75, -44, -52, 21, 56, 5, 64, -65, -48, -69, -52, -2, 49, 31, 21, -19, -53, 16, -36, -65, -19, -14, -28, 27, 13, 56, 12, -34, -63, -49, -75, -65, -20, -52, 32, -40, 27, 20, -32, 54, 24, -9, -26, -3, -56, 71, 51, -34, 9, -60, -26, 64, -1, 21, 15, -66, 0, -48, -27, 12, -24, -28, 20, 31, -5, -24, 64, -54, 69, -44, 73, 15, 20, -28, -63, 39, -35, 63, -73, 49, -75, -24, 35, -2, 70, -25, 7, -6, 0, 54, -70, 49, -50, 24, 2, 18, 73, -12, 38, 67, 19, 35, 6, -39, -69, 16, 75, -31, 2, -74, -57, 2, -23, 51, 73, -29, -50, 3, 41, 23, -19, 44, -4, 6, -8, 71, -52, -12, -17, 59, -21, 75, 19, 58, -40, 23, -3, -41, 68, 74, -42, -67, -2, 8, 59, -4, 53, -68, 74, 16, 30, -23, -18, -51, 56, 48, -56, -74, -40, 3, 61, 12, 2, 4, -6, 36, -51, 64, 68, -61, 62, -49, -53, -17, 32, -71, 54, 9, -66, 50, -51, 37, -51, 5, 61, -71, -23, -72, -70, 12, 4, 64, -52, -72, -10, 15, 39, 15, 4, 32, 27, -12, 56, 48, 46, 10, 52, 22, -56, 59, -6, -34, 20, 18, 46, 4, 20, -55, 7, 24, 32, -67, 12, 55, -64, -73, -5, 49, 15, 72, 3, -34, -16, -19, -62, -47, 66, 63, 50, -68, 46, -31, -28, -11, 60, -60, 68, 5, -39, -3, -47, 68, 5, 38, 46, 14, 38, -37, -15, -23, -41, 61, 17, 16, -34, 28, 44, -43, 16, 17, -38, -16, 61, 9, 48, 43, 25, 40, -30, 61, -41, -4, 53, 37, -41, 21, -26, 72, 59, 34, -28, -58, 20, 64, 32, 61, 14, 0, -60, -46, -59, -22, 12, 75, 60, -16, 41, 9, -53, -65, -6, -19, 7, -30, -59, 39, 64, -10, 35, 48, -52, -71, 63, 41, 68, 19, 27, 5, -58, 40, 34, -42, -60, -32, -44, -75, 28, 72, 9, 48, -69, -74, -49, 11, -31, -33, -26, -43, 32, -68, -73, 56, -64, 66, 21, -73, 7, -30, 7, 24, -67, -37, 58, -52, 7, -64, -52, -41, -68, 31, -71, -64, 32, -45, 21, 74, -2, 70, -47, -46, -74, -44, -68, -64, -56, 27, -62, 26, 70, 20, -27, -73, 58, -47, -49, -11, -36, -28, 21, -31, -73, 25, -20, 32, 54, 74, 30, -24, 69, 57, 3, 68, -65, 9, -72, -46, -40, -59, 53, -46, 34, -50, -45, 17, -22, -19, -72, 15, 28, 25, 59, 31, -28, -38, -15, -50, -40, -62, -1, -47, 70, -73, -56, -71, 9, -53, -44, 42, -38, -69, 69, 71, -45, -52, 12, 8, 4, 14, -54, -45, -39, -71, 59, 8, -34, -32, 32, 0, -19, -45, 28, -27, -45, 45, -23, 39, 68, 6, 3, -46, 13, -3, -51, 43, 20, 35, -27, -53, -27, -8, -23, 7, -3, -42, -61, 36, -1, 46, -40, 54, 75, 62, -49, -48, 31, 2, 67, 23, -68, -6, 50, 18, 64, 73, -17, 9, 32, 30, 31, -73, -54, -70, 9, 16, -39, 21, -23, 35, -10, 10, 13, -11, -4, 40, 16, -50, -36, 5, 46, -29, 73, 21, 65, 61, 18, -30, -8, -28, 75, -55, -28, -54, -50, 54, 37, -16, -1, -64, -56, 64, 22, 30, -25, -60, -8, 65, -35, 31, -8, -64, -73, -13, 30, 65, -29, -30, -43, 38, 17, -43, 59, 62, -24, -69, 40, -65, -9, -39, -55, 8, -52, 42, -40, -4, 55, 28, -15, -55, -17, 51, -46, -17, -38, 59, -30, 6, -47, 1, -31, 43, 33, -50, 27, -69, -46, -9, -61, 18, 25, -41, -52, 48, -75, -16, -31, 54, -64, 27, 74, -8, 0, -48, 49, 36, -67, -59, -34, -39, 17, 8, -74, -28, 31, 28, -24, 61, -59, -9, 1, 41, 25, 25, 12, 24, -67, 54, 2, -58, 3, -2, 7, -72, 25, -22, 37, 33, -5, -73, 67, -66, 9, 68, -18, -38, 18, 31, -55, 34, -54, 22, -3, 45, -31, -67, -7, -25, 62, 68, -8, -12, -10, 72, -9, -63, -25, -48, 43, 43, -48, 34, 52, 34, 24, -44, 72, -34, 63, -59, 73, -69, 36, -6, 51, -71, 1, -34, -21, -15, -42, 44, 48, 21, 41, -39, 33, -62, -14, 0, 56, 12, -44, 30, -30, 53, 62, -36, -59, 47, -21, -62, 53, -61, 6, 27, -56, -71, 68, -4, -11, -51, -35, -40, 45, -70, -6, 1, -59, 56, 74, 72, -8, -45, 26, 35, -70, 10, 73, -53, -21, -24, -40, -45, -10, 39, 57, 9, 43, 49, -72, -45, 73, -32, -12, 41, -29, 57, -34, -13, 35, -36, -19, -51, -8, -71, 60, -2, 15, 57, 20, 67, -43, 53, -54, 20, 15, -73, -48, -20, 50, -45, 10, 45, -2, 71, 10, 42, 53, 49, -47, 12, -62, 9, 37, 3, 11, 19, 74, -52, -2, 18, -60, 28, -6, -39, -28, -67, -38, -3, -12, -64, 27, 72, 56, -53, 67, -9, 64, 42, -38, -59, -23, -25, 23, -64, 52, -41, 28, 50, -18, -50, -9, -5, 51, 60, 32, -55, 66, 69, 18, -24, -73, -33, -30, 58, -10, -40, -29, -24, 75, 9, -7, -24, 57, -62, -13, 31, -30, -61, 6, 26, -38, 72, -55, -63, 54, 52, -44, 42, 43, 49, -60, 45, -62, -16, 26, 3, 19, 70, 55, 16, 1, -30, 68, -17, -19, -23, -62, 27, -10, 17, -23, 27, 11, -5, 38, -11, -30, 67, -47, -63, 40, -33, 56, 53, 26, 4, -21, -33, -4, -44, 58, 73, -1, 48, -22, 55, -50, -9, 4, 15, -69, 54, -36, 17, -26, 75, -71, 19, 66, -43, 29, 28, -3, 7, 4, -53, -67, 56, -13, 5, -64, -30, 2, 10, -58, 55, -13, -35, -32, 67, 55, -26, 43, -58, 65, -59, -61, 69, 33, -70, -52, -15, 33, 21, 67, -41, 41, 74, -61, -47, 3, -52, -2, -71, 33, 13, 57, -57, 54, -53, -68, 31, -3, 50, 46, -16, 65, 61, -23, 22, 66, -2, -69, 21, -59, 72, 54, 58, 70, 68, -67, -5, -59, 4, -3, 47, -59, -22, 65, 68, 0, 70, 24, 70, 45, -8, -24, 34, -23, 28, -20, -35, -51, -15, 60, -35, -21, 38, -55, -29, 28, -47, 41, 44, 32, -38, 14, 49, 13, 1, 39, -65, -4, -13, -70, -35, 53, -21, 72, -46, -70, -26, -5, -46, 34, -23, -8, -65, -61, 13, -19, 40, 39, -54, 7, -4, -19, -55, -33, 69, 21, -70, -71, -61, -9, -68, -23, -32, -14, -27, -5, -9, 23, 63, 18, -21, -36, -65, -10, -24, 23, 46, -59, -14, 66, 23, 55, -29, 43, -54, -35, -14, -50, -31, -1, 14, -26, 51, 57, 35, -51, -26, -51, 45, -38, 42, -52, 1, 52, 13, 53, -3, -18, 69, 57, -28, 14, 36, 18, -21, 56, 58, 40, -72, -51, -37, 17, -2, -63, -4, -44, -39, 45, -22, -70, -69, -56, -49, 6, 70, 40, -17, -9, -56, -26, -30, -9, 63, -71, -67, -36, 58, 65, -72, 61, -62, -35, 0, 10, -23, 71, 39, 11, 38, -59, 14, 43, -42, 40, -27, -48, 2, 29, 17, 21, -75, 62, -64, 63, 64, -57, -51, 46, -68, -50, 31, -57, -10, -47, 26, 40, -54, -13, -27, 60, 3, 62, 27, 35, 25, 73, 62, -51, 26, 1, 44, 26, -14, 55, 11, -26, 71, 35, -55, -75, 60, 49, -56, -27, -73, 43, -65, -52, -45, -16, -70, 31, -32, 30, -10, 66, 27, -25, -60, -25, 51, 59, 74, -39, 36, 9, 9, 30, -34, 27, 30, -51, 0, 47, -3, 0, 15, 5, 22, 45, 64, 25, 0, -45, -20, 64, -57, -71, -37, -42, -20, -64, -61, -22, -29, 49, 61, 55, 3, -49, 6, -45, -25, -72, -73, 45, 4, 17, -25, -52, -16, -39, 48, 57, -11, -50, 45, 8, -45, -70, 39, 8, -58, 54, 59, -12, 25, 44, -33, -48, 69, 48, -20, -34, 51, -18, -64, -23, 72, -16, 0, -20, 20, -29, -40, -66, -4, -71, 17, 26, -67, -20, -42, -50, -44, -58, 13, 56, 59, 53, -70, 52, 23, -14, -57, -4, 41, -48, 49, 38, 11, -29, -60, -47, 17, -25, -40, -62, -22, 50, 37, -14, -45, 69, 9, -16, -67, -54, -37, 67, 72, -32, 42, 19, 27, 58, -61, -9, -66, 61, -47, 18, -43, -34, 44, 47, 15, -71, 60, 68, 54, 20, -24, -69, 13, 60, -9, 21, -72, 29, 12, 75, 70, -22, 18, 20, -40, 30, -65, -33, 16, -39, 58, 48, 2, 27, 19, -59, 31, 2, -69, 9, -54, -18, 16, 34, -36, -71, -23, -33, 31, 64, -36, 23, -35, 55, -33, -2, 10, -25, 41, -52, 9, 23, 69, -64, -28, 10, -50, -73, -66, -45, 10, -45, 12, -52, 62, 50, -48, -37, -61, 56, -50, -23, 3, -12, -44, 44, 61, 39, -59, 24, 62, 26, -30, 53, 35, 17, -12, 60, 18, -3, -61, -48, 26, 25, -25, 10, -3, 0, 47, 11, -20, 72, 63, 58, -18, -58, 24, -33, 56, 41, 65, 41, -9, -43, 16, -52, 47, -72, -68, -11, -1, -55, 16, -53, 43, 66, 32, -36, -10, 3, 48, 43, -3, 34, 26, 54, 51, -28, -56, 29, -63, -69, -8, 1, -37, -67, 24, -66, -66, 30, -3, 6, 48, -63, 28, 15, -74, -15, 52, -11, 61, 24, -43, -17, -20, 56, -41, -47, -48, -22, 56, -37, -16, -28, 37, 20, -22, -16, 28, -14, -62, -51, 67, 59, -39, 18, -2, -40, -75, -28, 23, 61, 69, 55, -32, -26, 33, 1, 2, 58, 52, -20, -57, -41, 26, 56, 54, -72, -36, 6, -13, -25, 28, -23, -44, 63, 68, 27, -53, 68, 74, 45, 53, 67, 22, -56, -37, -21, 20, 39, -40, -4, -57, -22, 30, 44, -42, 7, 46, -5, -63, -45, 43, 39, 7, 72, 26, -1, 23, 48, -9, 21, 16, -33, 11, -40, -14, 49, 13, -70, 12, 48, -1, 29, -50, -48, -3, -18, 34, -35, 50, 44, -4, 16, 7, -73, 12, -43, 0, -40, -72, 64, 54, 17, -45, -11, 52, 16, -39, -13, 19, 46, -41, -59, -1, -17, -32, 70, 38, -74, -41, 10, 43, 30, -52, -25, 31, 34, 5, -47, 67, 8, -59, 45, -53, -30, -43, 73, 59, -9, -16, 1, -39, 17, 17, 34, 75, 58, 28, 35, 59, 60, -33, 26, 13, -9, 74, -34, -53, 4, -6, -62, -66, 8, 56, -43, 53, -65, -46, 35, 1, 13, -40, 38, -46, 52, -6, -49, 32, -54, 59, 15, -72, -49, -37, 16, 15, -40, 57, 37, 39, -27, 48, 48, 57, 28, -73, 32, 37, -44, -9, -38, 43, 24, 73, 70, -2, -9, -56, -46, 12, -73, 42, 14, -49, -70, -46, 41, -35, -66, 0, -74, -18, -30, 47, -39, 72, 50, 69, 33, -72, -18, 70, 44, -69, 68, 39, 4, -19, 56, 32, 67, 58, -2, 5, -68, 3, 34, 48, 41, 41, -29, 40, -52, 16, 12, -16, 10, -16, -25, -33, -15, 33, -40, -46, 37, -50, 66, -37, 6, 46, 70, -3, 26, -9, -74, 33, 67, 34, 4, 33, -1, 48, -5, 20, -14, -71, -71, 72, -12, -23, -37, 47, -68, -2, -75, 42, 21, 64, -70, -48, 32, 73, 22, -18, -12, 24, -62, -22, -20, 15, -67, 52, -13, 3, -3, 48, 8, -1, 44, 69, 51, -70, 40, 59, 1, 38, 25, -53, 26, 28, -28, -18, 24, 69, 38, -66, 17, 49, -13, 70, -12, -5, 47, 48, 74, -32, 20, 4, 42, -13, -3, 15, -10, -40, -2, 66, 73, -54, -65, 24, 49, -18, -72, -3, -24, 39, 7, 66, 10, 69, 61, 71, -13, 32, 43, -15, 73, -12, 64, 37, 48, -17, -24, -38, 18, 50, -50, 16, 69, -39, -38, 42, 18, -37, -38, 69, -75, 42, 58, 10, 33, 43, 6, -56, -3, -27, 2, -6, 34, -10, -45, 4, 47, 6, 41, -11, -22, 67, -71, -29, -50, -36, -64, 43, 3, -29, 35, 1, -63, 17, -65, 43, -18, 14, 63, 54, 61, -11, -28, 17, 53, 0, -54, 24, -72, 62, -63, -20, 51, -60, 24, 74, -21, 35, 40, 55, -72, -1, -20, -60, -62, -11, 59, -5, -75, 44, -29, 61, -43, 18, 3, -66, -60, 24, 31, -57, 8, 44, -2, -18, 59, -53, -20, -40, 55, -56, -62, 59, 16, -7, 72, 27, 55, 53, -54, 56, 21, -8, 41, 52, -68, -34, 59, -55, 63, 15, -36, -4, -17, 35, 51, -36, 55, -47, -3, 33, -29, 10, 16, 62, -72, 10, 14, 56, -12, 33, 36, -69, -52, 0, 58, -47, 39, 42, -26, 27, -21, 11, -55, 37, -32, 69, 74, -52, -54, -5, 56, -8, -70, -6, -23, -69, -74, 64, 62, -13, 19, 21, -6, 40, -55, -26, 69, 59, -62, -35, 8, -8, 49, 28, -49, -59, 21, -51, -36, 41, 18, -58, -43, 23, 9, 9, 29, 11, -3, 13, 73, -61, -42, -11, 54, -24, 39, 45, -42, 50, -66, 41, -33, 56, -8, -9, 73, -65, 16, -41, 51, -44, -25, -67, 54, 59, 15, 5, -6, -65, -60, -10, -51, -26, 54, -75, 23, 17, 46, 56, -10, 53, 20, 32, 34, -64, -55, 31, -54, 36, 63, 71, 65, -40, -74, 43, -56, 16, -30, 11, 24, -14, -75, 46, 33, 53, 47, -20, -8, 17, -41, 57, -6, 54, 13, -48, 63, 34, 56, -69, -8, 42, -74, -20, -74, -73, -53, -57, 17, -9, 30, -35, 50, 28, -64, 5, 5, 56, 60, 73, -3, -59, 54, 64, 70, -10, -59, 55, -54, 70, 62, 11, 34, 63, 66, 36, 66, -64, 54, 7, 2, 6, 45, -26, -41, 56, 54, 37, 34, 36, 34, -45, 53, 11, -56, 45, -75, -42, 25, -56, -48, 11, 30, 62, -2, 19, 20, -14, 30, -4, 66, -46, -73, 36, 3, -41, 14, -21, 71, -27, -61, 30, 1, 65, -37, 20, 35, -39, 51, -18, -20, -74, 68, -68, 61, -12, 26, 5, 48, -22, -75, 38, 5, -75, -2, -70, -41, -65, -16, -45, -17, -3, 58, 59, -14, -55, 2, -55, -21, -23, 2, 34, -22, -8, 39, -39, 56, -12, 41, 26, 41, 40, -12, -31, 40, 60, -26, 75, 70, 32, -48, -25, -47, -68, -44, 14, -50, 31, 33, 4, -69, -43, -38, -18, 25, 74, 19, 3, -14, -16, -47, -50, -52, 14, -6, 62, -2, 41, 59, -10, -3, -65, 38, 23, -58, 70, -40, -33, 23, 66, 46, 29, -53, -70, -64, 45, -72, 30, -30, -10, -64, -4, 13, -42, -65, -69, -56, 6, 45, -73, 70, -33, -65, 32, 63, -50, 24, -53, -10, -28, -63, -42, -75, -42, -37, -66, -73, -36, 37, -27, 27, 49, 44, -36, -69, 52, -32, -52, -17, -62, -50, -25, -22, -42, -69, -35, -17, 31, -14, 46, -75, -4, -72, 74, 29, -36, -69, 30, 1, 43, -75, -47, 16, 42, -10, 20, 17, 32, 43, 73, 45, 66, -28, -55, -52, -22, -17, 4, -69, 44, -26, -71, -37, -25, -72, 65, 14, -66, 19, -60, 52, 17, -34, -9, -18, 29, -65, 74, -15, 54, 71, -48, 44, -33, -30, 66, 18, 29, -6, 25, -3, 42, 29, 33, -59, 30, 23, 29, 39, -36, 42, 14, 57, -70, -73, -39, 34, -63, -41, -58, 66, -48, -33, 33, -6, 13, 23, -64, -34, -61, 34, 36, 54, -14, -6, 69, -60, -61, 22, 53, -22, -12, -11, -43, -7, -9, -7, -51, 3, 25, -36, -8, 52, 7, -51, -32, -56, 45, -22, -17, 57, -64, -59, 36, -3, 8, 29, 13, 22, -27, -12, 74, 36, 52, -45, -49, -33, 22, -27, 45, -29, 13, -39, -52, -56, -17, -9, -39, -48, 44, 17, -68, 54, 31, 43, -25, -36, -4, 61, 59, 42, -27, 57, 0, -51, -65, 26, -9, 32, 72, -41, -73, 9, -5, -52, 26, 52, 13, 60, -74, -21, -1, -67, -43, -45, 49, 6, -8, -31, -11, -25, -65, 38, -45, 10, 60, -37, -42, -26, 68, -47, 8, 70, 35, -75, -59, -16, 52, 27, -32, 52, -70, 43, 60, -39, 71, 34, 42, -13, -75, -47, 35, -66, 64, 63, 17, 49, -50, 49, -53, -58, 75, 28, -65, 34, 28, -51, -58, 3, 51, -16, -21, 56, -51, -39, -61, -56, 68, 54, 4, 67, -68, -37, 74, 71, -49, 13, 44, -26, -14, 64, -10, -17, 16, 0, -58, -33, 24, -43, 45, -1, 14, -54, -23, 38, -20, -8, 55, -29, -30, -19, -38, -23, 20, -42, -29, 44, 46, -61, -60, -45, -74, 5, 13, 15, -71, 30, 57, 26, 61, 24, -53, -1, 43, -2, -40, -52, 65, -63, -8, -43, -6, 29, 8, -64, 62, 54, 53, 32, 66, 68, 62, 65, -2, -2, 5, 0, -50, -14, -51, -65, -67, -31, 8, 51, 42, 43, 72, 29, 55, -12, 62, -29, -61, -8, -18, -75, -30, -41, 31, -42, -50, 15, -52, 21, -63, 28, -57, -39, -64, -33, -29, -56, 12, 54, 69, -24, 19, 65, -70, -3, -22, 65, 43, -8, -19, -52, -9, 24, -20, -56, 55, 5, 32, -73, -50, 43, 28, -33, -72, 38, 9, -26, 57, -57, -49, 50, -7, 45, 38, -2, -36, -60, -13, -68, 5, 41, -45, 69, -13, 8, -65, -34, -62, 43, -33, -39, 10, 70, 3, 11, 32, -65, 58, 12, -49, -67, -16, 19, 52, -54, -61, -60, -41, -1, -55, 38, -36, -27, 31, 26, 57, 42, 66, 68, 7, -43, -49, -61, -51, 30, 25, 55, 38, 7, -9, 62, 14, 50, 6, -10, 70, 20, 3, -47, -56, 24, 66, -19, 72, 20, -70, 51, -16, 71, 43, 66, -48, 70, -73, -24, 22, 25, -47, -16, -44, 19, -30, 45, -8, 49, -43, -16, -8, 36, 12, 9, -18, 1, 65, -22, -57, 70, -46, 2, 65, 70, -10, -61, 64, -8, -11, 10, -59, 17, 67, -30, -39, -40, -62, 26, -69, -32, -66, -2, -74, 19, -69, -17, -56, 70, 35, -38, 64, 62, 37, 52, 56, -49, 66, 45, 16, -21, -23, 30, 72, -33, -75, -45, 2, -64, 54, 8, -21, 63, -71, -19, 4, -67, 39, 24, -73, -2, 59, 67, -16, 21, 41, -35, 45, 31, -68, -16, -67, -18, -62, -73, 24, -62, -43, -50, -53, -67, 32, 2, 71, 34, 58, -1, 42, 19, -55, 43, -58, -73, 32, -1, 21, -3, 37, -12, -48, 42, 47, -42, -51, 61, -40, 48, 72, -10, 72, -56, -2, 26, 21, -9, -16, 1, 64, -52, -56, -67, 66, -41, -67, 22, 32, 27, -59, -9, -60, -31, -42, 62, 0, -18, 45, 36, -48, 42, -50, -52, 61, 24, 49, 4, -61, -45, -71, -73, -23, -54, -66, -35, -21, -60, 61, -65, 43, -74, 1, 58, -32, 34, 42, 44, -62, 12, 4, -34, -22, 27, -13, -39, -25, -39, 38, -12, -11, 42, -12, 39, 61, -5, -71, -36, 11, 63, -26, -22, 64, 49, -42, -45, 5, 75, 74, 19, 9, 0, 60, 60, -49, -29, -55, 0, 5, 58, 61, 68, 22, -27, 31, 8, 44, 33, 45, -23, 20, -58, 30, 7, 66, 61, 37, -5, 58, 35, -64, -8, -43, 69, -24, -17, -37, -5, 56, 43, -25, 41, 33, 73, -63, -13, 3, 54, -58, -30, -45, 38, -13, 60, -33, -23, 43, -72, 46, 25, 36, 57, -59, 68, 51, -9, -27, -62, 61, -48, 54, -40, 68, 10, -45, -73, 72, 31, 56, -62, -74, -65, 49, -12, 68, -62, 39, 35, -59, 9, -15, 50, -10, -1, 42, -37, 65, -62, -24, 50, -35, -47, -67, -45, 38, -37, -42, 34, 68, -64, 45, 69, -53, 17, -19, -63, 30, -56, 46, 47, 26, -45, 19, -59, 29, -16, -23, 19, -3, 29, -9, 35, 57, -1, 65, 19, 36, -55, -25, 28, -43, -58, 21, -23, 34, 75, -13, -11, -58, -43, -42, 41, -15, 52, 57, -61, -40, -41, 31, 30, 61, -56, -13, 40, 19, -25, -19, -23, -5, 31, -71, 25, 48, 23, 75, 7, 20, -15, 69, 37, 17, -51, 3, -73, -75, -18, -61, -41, 14, 43, 62, -3, 62, -26, -39, 3, 24, 17, 55, -59, -30, 59, 40, -59, 6, 39, 21, -49, -52, 14, 61, 39, 38, -14, 39, 36, 42, 53, 68, -20, 18, 55, 51, 4, -49, -64, -70, 50, 27, 60, 64, 70, 42, 28, -65, -28, -10, 31, -4, 11, -33, -20, -26, -71, 39, -65, 39, 5, 63, 31, 59, 3, 10, 34, -68, 34, 43, -63, 8, -8, 70, -3, -13, 36, -53, -3, -69, 12, -49, 0, -54, -7, 55, -5, -4, 17, 6, -41, -54, -9, 65, -71, 70, -2, 36, 75, -44, 4, -66, 38, 71, -72, -43, -18, 40, -21, 53, 44, 65, -72, -32, -65, -4, -54, 3, 67, 38, -67, -52, 59, -2, -62, 62, -10, 9, 22, -11, 40, -52, -4, 0, -58, -3, 32, -1, -39, -64, -26, -71, -75, -23, -29, -65, 47, -8, 11, 36, -46, 20, 60, -63, -60, 71, 72, 3, 4, 19, 67, -34, 40, -15, 42, 57, 57, -2, -21, -59, 7, 28, -57, 7, -72, -11, 15, 48, 56, -49, 8, -66, 44, -10, -55, 57, -15, -59, -16, 62, 33, -27, -47, -2, 33, 70, -21, 12, -8, 33, 28, 75, -16, 47, 4, -13, -42, -58, -41, -61, -34, 40, -54, -68, -45, -34, 64, 13, -17, -28, 0, -62, 18, 28, 11, -27, 20, 64, 60, -66, 21, 13, -69, -73, -18, 11, -11, 15, 26, 21, 27, 67, -16, 49, 74, 14, -61, 60, -51, -5, -46, 24, 9, 47, -26, -58, -56, 67, -70, -74, -74, 25, 12, -68, 27, 69, 16, -61, 7, -34, 33, -42, -45, -59, -69, -49, 28, -54, -65, 53, 14, -38, -1, -55, -67, 47, -37, -50, 38, -32, -50, 39, 66, 37, 45, 16, 29, -15, 28, -40, 27, -15, -7, 55, 2, -2, -69, -46, 17, -59, -71, -45, -21, 4, -24, -15, -27, 12, 9, -65, 53, 34, 48, 44, -7, 17, -18, -54, 75, -66, -19, 24, -6, 48, 4, 71, -30, 10, -52, 60, 24, -48, -63, -75, 29, -12, -16, -74, 73, 68, -63, 51, 24, 58, 17, -59, -3, 74, -37, -4, -68, 17, -55, 1, -11, 24, -5, 32, -44, 18, 14, 55, 43, 27, 56, -3, -63, -36, -2, -65, -46, 8, 61, 53, -10, 2, 67, 60, -2, -48, -19, 5, 45, -1, -72, -44, -53, -2, 62, -22, -62, 0, -45, 57, -51, -65, -24, -38, -28, 49, -30, 1, -18, -45, -24, 45, 30, -32, 30, -48, -7, -67, 32, -38, 7, 33, -8, 27, -46, -24, -73, -33, 49, -43, -54, 74, -34, -3, -42, 11, -31, 3, -63, 24, 33, -14, -7, -15, 27, -55, 12, -55, -49, -34, -20, 33, 72, 45, -18, -50, -55, -16, -9, 68, 15, 12, 66, 56, -68, -52, -11, -24, 26, -1, 75, -19, 61, -10, 39, 10, 11, -27, 30, 35, 12, -67, -7, 8, 51, 50, 34, 72, -43, -51, 64, 47, 34, 52, 25, 41, 73, -62, -61, 21, 13, -64, 75, -4, 2, 38, -70, -65, -65, 34, 45, 22, 40, -40, -48, 15, -67, 61, 9, -35, -68, -5, -66, 40, -31, 34, 3, -34, 45, 18, 62, -20, 27, 61, 49, -47, 21, 55, -39, 29, 11, -69, -25, -27, -36, 1, 63, -28, -16, -5, 10, -8, 65, 19, -44, -41, -25, 32, -2, -57, -26, -15, -2, -74, -32, -30, -48, 65, -53, -11, 18, 33, -7, 67, -70, 32, -8, 66, -71, 51, -15, 12, -35, -27, -44, -6, 5, 6, -49, -73, 22, -2, -13, -55, -3, 29, -10, 25, 18, 12, -64, -42, -33, 4, -53, -30, -42, 14, -42, -40, -12, 17, 48, 26, 65, -72, -55, -8, 7, -31, -6, -46, 42, 55, -28, -36, 8, 35, 62, -52, -31, 71, -21, 9, -1, 2, 52, 30, -62, -66, 66, 1, 26, 38, -50, 13, 39, -30, -71, -32, 14, -1, -5, -22, -24, 40, 15, 59, -3, -1, -71, 41, -6, -17, -28, 66, 60, -52, 21, 74, -42, 11, -3, 57, -29, 22, -5, -66, 65, -1, -25, 1, 71, 46, 55, -29, 10, -8, -48, -68, 67, -44, 46, -15, 13, -59, -24, -5, -36, 70, -7, -5, 5, 64, -23, 49, 8, 47, 56, -2, -32, -45, 74, -36, 74, 51, 10, 7, -32, 38, 14, -43, 67, -18, 17, 4, -2, 66, 75, 36, 60, -10, -45, -13, -22, 7, -40, 62, -24, -62, -18, 20, -31, -20, 59, -33, -46, -9, 49, -3, -49, -15, 29, -57, 41, -32, 20, -39, -43, 19, 72, -61, -68, -50, 0, -17, 30, 33, -33, -69, 47, 24, 24, -62, -73, 5, -20, -44, 71, -48, 26, -53, 10, -23, -37, -27, 18, 58, 10, 48, 0, 4, 63, 5, 29, -15, 63, -16, -58, -47, -12, 62, 50, -66, 75, 52, 14, -22, -70, 7, 5, 29, 27, -63, -72, 65, -14, 20, 46, 71, -8, -32, -1, -23, 48, -49, 37, 33, 8, 53, 61, 69, 39, 36, -73, 39, 10, 14, -59, 16, -55, 19, -33, 48, 31, -29, 35, -61, 64, 5, -66, -20, 48, 7, 31, 18, 31, -8, -24, -37, -33, -39, -44, -69, 70, -44, 43, 5, 45, 57, -57, 63, 0, -15, 33, -47, 29, -7, -32, 17, 73, -25, 71, 44, 57, 26, -14, 12, -60, 35, 48, -17, 72, -74, -11, 64, -43, -46, -7, 75, -65, 11, 61, 10, 70, 18, 36, 23, -65, -72, -37, -69, -21, -42, 48, -42, 57, -42, 46, 72, 67, 16, -21, 61, 18, 41, 49, 48, 68, -33, 46, -73, 51, 31, 10, 45, -27, -29, -9, -18, -26, 29, -14, 26, 60, -42, 60, 41, -11, 28, 37, -20, -32, -61, -35, 59, 53, -61, 32, 46, -21, 2, 48, -46, -45, -19, 73, 1, 27, -12, 58, 74, -59, -32, 25, -75, -1, 7, 39, 64, -41, 0, -32, 0, 12, 7, -16, -10, 19, -60, -42, 71, 15, -72, -51, 45, -16, -54, -30, -65, 7, -49, -66, 23, -8, 32, 21, 67, -37, -16, 53, -5, 58, -57, 68, -6, 25, -24, 57, -34, -11, -63, -39, -74, -59, -16, 44, 0, 3, -63, 9, -65, -37, 16, 33, 28, -30, -23, 19, 8, 36, -4, -75, 16, 15, 68, -67, -38, -33, 65, 4, 29, -75, 38, 31, -59, -54, -1, 14, 25, 11, -55, 35, 47, 36, -10, 0, -70, 40, -59, 11, 1, 13, 9, -61, -50, 0, -53, -15, 42, -63, 62, -5, -65, 25, -50, -51, 46, 23, 38, -7, -42, 57, -50, -72, 15, 14, 3, 21, -22, 19, -46, 52, -46, 39, 67, -23, -37, -62, 38, -73, -52, 24, -3, -42, -29, 21, -18, -60, -34, -57, 8, -3, 75, 34, 0, 14, -28, -73, -43, 23, 20, -15, 0, 49, -52, -9, -49, -16, 4, 62, -16, 28, 8, 54, 61, 53, -1, -32, 68, 38, -14, 0, -40, -17, -44, 33, 72, 1, 34, -48, -51, -22, 12, 24, -51, 33, -61, -27, -59, 16, -41, -2, -32, 41, -24, -46, 18, 51, -5, 10, 11, 54, -68, 44, -41, -38, 2, -47, 38, -40, -20, 60, 11, 67, 6, 35, 24, 20, -67, 38, -39, -35, -40, 2, -72, 10, 29, 21, -17, -52, -47, 69, 75, -41, 38, -42, -4, -36, -13, -44, -3, 42, -59, -68, 32, 22, 42, -22, -35, 48, -61, -1, -64, -28, -75, -61, 57, 30, 34, -36, 51, 62, -42, 49, -57, 69, -69, 14, -43, -9, 46, 27, -44, 60, 34, 63, 4, -2, -37, 44, -29, -25, -35, -18, 23, -36, -6, 2, 67, -48, 42, 42, -63, 73, 15, -45, 66, 20, 45, -55, -65, 13, 45, -34, -5, 3, -49, 74, -75, -12, 41, -31, 38, -70, 24, -15, -33, -57, 63, -42, -30, 27, -75, -20, 22, 13, 11, 10, -45, -22, 28, -34, 66, -3, 5, -17, 75, 30, -19, 73, -58, -56, -35, 55, -52, 64, -37, -10, -71, -52, 24, -27, 50, 22, 28, -6, -43, -37, -72, -12, 16, 31, 27, 4, -48, -46, 62, -51, 59, -34, -56, -75, -17, -18, 54, 6, -29, -59, 72, -27, -36, 18, 21, -62, -38, -26, 5, -6, 10, 8, 55, -51, -37, 6, 28, -12, 36, 13, 10, 17, 52, 27, 18, -41, -66, -6, 41, -22, 10, 35, 26, 49, -25, -28, 60, 12, 19, -11, -72, -49, 72, 59, -25, -43, -13, -74, 18, -55, 12, -48, 38, -14, 52, -22, 20, 61, 47, -17, -37, -19, -60, 65, -48, -10, -41, -66, 75, 51, -2, -72, 75, -8, 60, -27, 22, -31, -26, -36, -10, 59, -11, -50, -31, -35, 3, 62, -49, -28, -30, -13, 26, -17, -24, 53, 47, 8, 62, 46, -17, -18, 47, -19, 47, 29, 29, -7, 74, -75, 30, -12, 59, -57, 13, -50, -19, -62, -64, 5, -15, -21, 68, -67, 38, -34, 59, 9, 50, 45, -23, -45, -51, -51, 11, 71, 53, -36, -12, 49, -36, -60, -39, -55, -42, 47, -30, 12, 58, -20, -58, -33, 34, -68, -27, -6, -27, -44, -73, -55, 74, -20, -24, -53, 2, 62, -58, -23, -51, 3, -49, -12, 18, -15, 7, 49, -43, 52, -16, -63, -46, -1, -20, 64, 6, 26, -18, 52, 58, -17, 73, 56, 36, -27, -72, -40, -43, -57, 12, -21, 20, 36, 41, -40, -54, -28, -68, -24, -54, -9, -12, -24, 63, 41, -36, -7, -8, 19, -33, -28, 75, -36, -48, 33, 10, -47, 68, 41, -30, 3, -56, 63, -37, 60, -55, -18, -46, -48, 33, -24, 16, -56, 27, 3, 58, 64, 69, -28, 5, -39, 19, 3, 0, 45, -40, -65, 71, -47, 49, -35, 31, 68, -50, 69, 51, -29, -26, -71, -2, -69, -22, -63, -52, -73, 15, -69, 64, 9, -24, -6, 45, 71, 70, -33, 40, -46, -25, 35, -18, -52, 74, -65, -61, -52, -73, 65, -6, -24, 67, 66, -20, -32, -73, 4, -30, 15, 8, -41, -52, 59, 26, 66, 52, 20, -44, 14, 47, 4, -28, -48, 28, -30, -38, 40, -9, -36, 27, 59, 15, 16, 49, 71, 59, 49, -3, -48, -12, -71, -14, 10, 61, -66, -2, 38, 27, 29, -24, -4, -42, 23, 23, 59, 66, 61, 21, -18, -51, -28, -35, 38, 63, -64, 33, 47, 60, -46, 74, -30, -44, -18, 55, -59, -11, -22, 52, -62, -71, -47, 9, -40, 49, -43, -59, 40, -60, 37, -54, -36, -67, -16, 75, 70, -5, 32, 39, -23, 59, 35, 22, -63, -59, 0, -48, 3, 53, -72, 14, 55, -46, -53, -62, -72, -23, -46, 43, -8, 67, 62, 30, 73, -30, 29, 67, 38, -16, 30, -61, -35, -11, 34, -22, 3, -42, 5, -72, -67, 6, 17, 62, 36, 38, 75, 39, -61, -47, 4, 5, -58, -10, -41, -60, 33, 61, -69, -5, -31, 35, 7, 10, -52, -35, 61, 25, -3, -12, 28, 5, 69, -30, -9, 27, -68, -12, -12, -56, 17, 67, 22, 34, -21, 54, 49, -64, 40, 54, 4, -69, 13, -67, 14, 34, -28, -1, -17, 44, 62, -64, -29, 56, -21, 36, 5, -16, -52, 69, 1, 38, 60, -52, -3, -38, -74, -32, -29, 39, -56, 49, 46, 30, 57, -16, -11, -47, 59, 45, 70, 43, 56, -34, 21, -43, 75, -49, 16, -53, -56, -58, 59, -74, -37, -22, -37, -36, 19, 8, -74, 39, -19, 47, -7, -38, -47, 55, -11, -64, 25, -17, 53, 3, 22, -2, 36, 21, 22, -26, 42, 41, -11, 23, 41, 27, -75, -74, 65, 19, 9, 66, -18, 65, 35, 49, -50, 63, 28, 12, 73, -25, 68, 50, 54, 15, -30, 14, -42, 68, 61, 73, 31, -25, 20, -4, 75, 20, -2, 62, -38, -71, 52, 19, 68, 11, -10, -60, -1, -59, 27, -4, -9, 17, -32, -31, -46, 13, 56, -12, 5, 42, -17, -39, -61, -74, 30, -62, 19, -50, -75, 56, -45, 50, -2, -55, -16, 63, -40, 56, -72, 60, -26, -7, 1, 17, 37, 31, -48, 16, -59, 33, -18, -1, 67, -6, 0, 19, 7, -56, 45, 5, 75, 73, -22, -5, -58, 37, -17, -23, 17, -16, -41, 66, 52, 35, 5, 12, -10, 32, -48, 6, -11, 7, -72, -22, -75, 3, 71, 5, 20, 40, -67, 18, 35, -14, -63, 52, -55, -7, -49, 37, 53, -15, 25, 27, -58, -46, -39, 8, 61, -14, -64, -27, 68, -61, 26, 66, 16, 21, -6, -42, -17, 0, 51, -58, 59, 62, 67, -72, -21, -60, 40, -46, 0, -11, 57, 16, 16, -60, -52, 1, 2, -43, 49, -6, -28, -2, -17, 61, -59, 50, -57, 0, -26, 68, 15, -43, 54, 7, -42, -43, 22, 71, -13, -55, -18, -34, 36, 73, -19, 57, -2, 58, -62, -30, -25, -17, 43, 33, -34, 59, 5, -17, -19, 54, -25, 72, -67, -47, 1, -34, -15, -55, -41, 45, -37, 16, -65, 72, 13, -8, 53, -67, -28, 65, -22, 22, -30, -57, -23, 10, -75, 57, 68, -19, 33, -33, -25, 39, -5, 49, -73, 53, 68, -39, 23, -45, 52, 31, -48, -13, -55, -73, -4, -7, 65, 47, -63, -42, 66, -12, 41, 66, -33, 33, -31, -75, 73, 18, 37, -8, -9, 40, -33, -19, 74, 63, 12, 49, 19, 37, -40, 39, 37, 29, -46, 25, 1, -33, 58, -11, 30, 23, -21, 70, -22, 21, 70, -25, -37, 32, 40, 28, -6, -69, -67, -8, 68, 18, -37, 11, -21, -1, -28, -59, -48, 2, 39, 26, 42, 21, -61, -6, -34, -9, -12, 19, -63, -19, 67, -27, -65, 31, -75, 4, 35, -68, 69, 27, 25, -43, -38, -73, 29, 8, -59, 54, -66, 55, 5, 49, 0, 17, -33, 39, -67, 28, -18, -57, -67, -27, -9, -57, -74, -10, 20, 36, -5, 12, -12, -56, 42, 23, -54, -7, -47, -38, -29, -40, -59, 49, -67, 14, -9, -27, -23, -3, -74, 32, 15, -68, -73, -72, -51, -74, -9, 42, 38, 61, -22, -52, -72, -58, 44, -51, 10, 73, -15, 55, -43, -1, 28, -34, -64, -57, 12, -14, 13, 11, -59, -48, 19, -59, -46, 41, -57, 20, 7, 56, 4, 59, -72, 7, -75, 45, 29, 9, 42, -62, -12, 75, 11, -60, -37, 22, -43, 50, -70, 45, -14, -54, 71, -71, -37, -51, 45, -19, 42, -26, -41, -30, -43, -40, 52, -44, -71, 4, 38, 47, 15, -50, 46, -50, -37, -67, 45, -7, 56, 51, -39, -34, 70, -44, -30, -43, -22, -63, 11, -58, -15, 45, -12, 15, -73, -38, 46, -68, 41, 6, 54, -19, 29, 22, 4, 68, 28, -28, -17, 8, -55, 19, 48, -61, 48, -60, -30, -52, -49, 56, -34, 11, 24, 27, -50, 26, 62, 70, 31, 28, 0, 9, -69, -46, -47, 8, -56, 54, 55, 0, -15, 75, -56, -43, -63, 67, -28, -18, -60, -2, -40, -21, -69, 57, -70, -43, 8, 67, -51, -37, 17, 24, 46, 21, 51, 72, -46, 68, 49, -69, -7, -42, -69, 10, -12, -57, 1, 33, -2, 14, -46, 33, 66, -40, 15, 71, -8, -55, 63, 14, -19, 2, -37, -51, -52, -64, -56, -25, -73, 68, -19, -5, -52, -15, -71, 9, 1, 3, -34, 74, -60, -7, 30, -70, 29, -33, -74, -57, -15, 62, 33, 39, -14, 69, 64, 9, -71, -70, 57, -71, 71, -37, -1, -57, 21, 1, 25, -55, -71, 64, -57, -58, -18, 46, -53, -67, -65, -54, -49, -5, -70, 57, -41, -8, 50, -55, -75, 53, -50, 56, 57, -55, -59, -21, -39, 37, 55, 59, 57, 57, 47, 74, 74, -49, 42, -56, -41, 53, -35, -16, -30, -29, -35, 2, 38, -62, 22, 36, 66, 45, 16, 45, 63, 32, -54, -52, -8, -74, -71, -29, 56, 52, -33, 55, -75, -66, 74, -42, 60, -39, 17, -48, 7, 55, 30, -33, 68, -24, -72, 56, -56, 17, 24, -69, -28, 45, -47, 37, 46, -43, -68, 25, -69, -27, 4, -68, -18, 0, -35, -36, 36, 55, -9, -34, 34, -57, 8, 25, -7, 9, 5, 12, -51, -47, 18, -4, 74, 46, -45, 42, -74, -38, -9, -68, 8, 68, -63, 63, -10, -23, -49, -51, -46, 16, -10, 64, 34, 71, 13, -49, 3, -60, 38, 25, -31, -21, -57, -35, -53, -27, -71, -52, 8, -6, -46, -59, -16, -34, -72, 50, 17, -45, 74, 46, 44, -14, 32, 2, -21, -31, 27, 57, -15, -13, 6, 27, 39, 22, 65, 62, 70, 67, -68, 3, -15, -41, 19, 45, -1, 22, 17, -60, 50, 15, 59, 16, 74, 16, -59, -23, 58, 43, -43, -35, -48, 36, 67, 67, -17, 54, 51, -23, 46, 56, 55, -47, -60, -4, 71, 14, -59, 12, 27, 64, -51, 10, 5, -53, -52, 21, 0, -69, -14, 32, -29, 11, -8, -39, 2, 50, -61, -25, -50, 58, -44, -73, -64, -31, -1, -69, 56, 15, 17, 7, 1, 41, -61, -70, 64, -37, 24, -14, -33, -68, -58, 13, 19, 7, 47, -55, -20, 62, -6, 5, 42, 25, 7, 51, 67, -72, 58, 47, 16, -3, -24, -58, -38, -10, -55, -50, 26, 45, 11, 68, 50, 26, 6, -7, -44, -25, 12, 11, -39, -70, -62, -74, 28, 18, 52, 19, 22, 32, -12, -38, -47, 39, -21, -9, -49, -2, 14, 53, -35, -52, 43, -61, 47, -29, 8, -75, 22, -56, 11, 56, -53, 22, 57, 50, -35, 34, -9, 62, -12, 52, -54, 17, 15, 1, -70, 39, 72, 17, 14, -39, 38, -18, -25, 8, 28, 58, 8, -28, 75, -56, -47, -54, 39, -68, 69, -72, 39, -18, 63, -48, -42, -66, 42, 46, 8, 45, 10, 4, -14, -52, 40, -53, 3, -61, 30, -46, 71, -38, 1, 68, -21, 27, -61, -57, 35, -70, -56, -2, -12, -68, 25, 21, -59, -11, -8, 24, -42, 75, -50, 20, -55, 65, 40, 24, -74, -6, 51, 70, 31, -24, 63, -67, -74, 75, -49, 36, -71, -30, -42, -10, -23, 57, -64, -9, -30, 1, -63, 4, -2, -38, -54, 18, -51, 61, -36, -49, -23, -61, -57, -70, -11, -70, -62, -10, -71, -36, -52, -68, 8, -19, -3, 58, -40, 6, -28, 4, -71, -16, -68, 2, 22, -49, -57, 44, -66, -18, 68, -14, -3, -64, -9, 61, -61, 5, -27, -58, 42, -4, -51, -28, 50, 19, -45, -65, -52, 2, 12, -50, 61, 17, 26, 5, 43, 44, -26, 50, -50, -36, -40, 20, -25, 24, 3, -10, -49, 51, 7, 67, -31, 29, -37, -56, -30, -7, -48, -7, 68, 39, 19, 52, -20, -31, -21, -55, -65, 26, 70, -40, 66, -48, 54, -35, 49, -19, 28, -75, -45, -43, 67, -1, 61, -48, 16, -46, 21, 43, 22, 11, 4, -37, -13, 57, 5, 42, -74, 15, -10, 69, 49, -20, -55, 27, 19, 68, -70, -29, 68, -42, 4, 57, 33, -13, -67, -29, 16, 27, -63, -39, -37, 16, -3, 23, -2, -73, -13, -3, 17, 53, -9, -12, -43, 9, -63, 51, -1, -57, -55, -9, -24, 22, -30, -69, -69, -23, -24, 23, -74, -12, 57, -36, -74, -22, 61, -1, -22, -30, 70, 69, -53, -17, -19, -22, 65, -6, -49, -11, 10, -29, 53, 61, 66, -52, 66, 73, -2, -34, 18, -1, 29, -1, 37, 28, 50, 20, -50, -47, 65, -56, -56, -63, 0, 0, -12, -11, 69, 14, 53, 3, 59, 29, -13, 49, 50, -25, 46, -28, 16, -12, 44, -33, 60, 5, 70, 33, -51, -56, 59, -61, -39, -73, -51, 36, 2, 10, -52, -6, -52, -75, 70, -71, 27, -21, 52, 1, 29, 20, 46, -33, -69, 15, 9, 64, -56, 2, 21, -31, 19, 4, -19, 56, 6, 5, 14, -69, -61, 37, 0, -40, 36, -8, -37, -13, 47, -61, 62, 0, 32, 32, 43, 38, -29, -26, 27, -9, 49, -28, 33, -7, 50, -64, -29, -20, 14, 58, -16, 26, 20, 59, 59, -22, -26, -54, 38, -55, -42, 24, 20, 66, -19, -15, 26, 25, 33, -25, -62, 6, 21, 46, 72, -5, 55, -35, 48, -7, -54, -43, -57, 39, -62, -73, -59, -13, -54, 54, 7, -20, 3, -50, -32, 57, 8, 67, 6, -35, -33, 20, 45, 63, -12, 39, -18, -32, -73, -48, 36, -52, -16, 53, 62, -2, 55, -73, 58, 74, 54, -10, -22, -19, 13, 19, -38, -55, 11, 42, -16, 51, -14, -49, 38, 49, 65, -58, -59, 67, -31, 51, -63, 29, 28, 74, -51, 5, 74, -69, 3, 53, -6, 55, -44, -71, -2, -8, -52, -69, -42, 7, 57, 19, 33, 17, -8, 20, 34, 7, 10, -72, -18, 22, 30, -66, 19, 52, 14, 15, 56, -59, -10, -27, 71, 22, -23, -8, -64, 0, -2, -31, -71, -22, 61, 37, 70, -25, -20, 27, 57, 65, 28, -37, 9, -18, -30, -50, -44, 59, 41, -64, 74, -45, -18, 69, 50, 35, -17, 61, -43, 57, -48, -38, -43, -63, 72, -51, -12, -24, 51, -31, -37, 3, 6, 46, 58, 51, 71, -64, 35, 34, -52, 33, 63, 3, 24, 37, -38, -68, 21, -5, 62, 48, 32, -59, 61, 28, -35, -27, -73, -61, 15, -35, 15, -55, -65, -2, 72, -71, 9, 29, 38, 30, -16, 25, -42, -68, -15, -7, -63, -70, 61, 72, 51, 17, -63, 36, -32, -24, -69, -32, -10, 22, 8, -71, 40, 17, 0, 34, 21, -68, -13, -19, 35, 46, -69, 68, 52, -11, -16, 62, -8, -31, 59, -33, 60, 69, -74, -50, -31, -70, -7, 32, 25, -75, 37, -10, 17, -41, -52, -40, -34, 9, 17, -74, -23, 21, 67, -47, -68, -25, -62, -1, 18, 72, 39, 2, 63, 38, 25, -43, 44, -58, 64, -7, -60, 23, 56, 33, 58, -73, 66, -52, 11, 7, -53, 63, -50, -61, -61, -43, -13, -50, 31, -71, -54, -7, 4, -69, -45, -47, -39, 72, -32, -50, -12, -16, 46, -32, -61, 26, -32, -71, 48, 52, 10, 70, 38, 35, -69, 52, 68, -6, -74, 21, -4, -55, -64, 74, -51, -35, -51, -14, -39, -7, 9, 24, 52, -21, 66, 66, -70, -44, 68, 53, -67, 2, 45, 46, -40, 52, 20, -48, -32, 19, 46, 37, 37, 58, 33, 61, -53, 58, -29, -19, -27, 55, -72, -53, -41, 69, -63, -38, -53, -73, -63, -45, 5, 57, -75, 40, 31, 20, 65, 74, -39, 35, 36, 73, 15, -9, 59, 35, -27, -46, -59, 19, -68, -58, 41, -36, -65, 53, 1, -43, 54, 11, -14, -17, -8, -14, -55, -52, -71, -66, -56, -37, 42, 53, -39, -20, -31, -56, -63, 17, -29, -49, -41, -22, -32, 75, 15, -22, 51, -60, 9, 29, 24, 68, -66, -59, -22, -46, -38, -20, -39, -19, 19, -75, -41, 53, -22, 3, 70, -9, -58, -35, 17, -24, 17, 61, -24, -44, -39, -51, -30, 43, 53, 69, 35, 62, -68, -64, -60, -33, -9, -26, 24, -68, -26, 56, 60, 28, -19, 54, -59, -4, -58, 33, 46, 32, 18, -56, 63, 53, -32, -45, 20, -55, -53, -20, -71, -48, -9, -56, -5, 55, -9, -59, 63, 38, 70, 45, -12, -25, 24, 4, 44, 39, -40, 14, -5, 53, 33, -20, 28, -75, 11, -27, -57, 31, 28, -53, 58, -59, -36, -25, 71, 30, -11, 58, -7, -17, 28, 54, 31, -26, -17, 0, -65, 18, -62, 5, -7, 45, 60, -54, 45, -7, -8, 62, -52, -56, -67, -71, -40, -27, -23, -47, -75, 42, -64, -9, -53, 37, -30, 54, -67, 26, -24, -57, -34, -13, 23, 32, -44, 5, 51, 75, 74, -33, 59, -56, -16, 67, -54, 17, -38, -1, 46, -37, -37, 55, 27, -15, 14, 70, -39, 22, 20, 10, 38, 59, 71, -15, 16, -49, 63, -9, -52, 61, 32, -69, -72, -62, 72, -51, 31, -42, 21, -1, -6, 59, -22, -54, -33, 67, -60, 1, 11, 34, -66, -27, 17, -71, 31, -45, -47, 18, 20, -23, 2, -24, -19, 5, -11, -23, 27, -58, 9, -27, 16, -75, -46, 67, -54, -6, 58, -40, 71, -9, 67, -71, 39, 6, -69, -8, 37, -41, -65, -19, 9, 10, 32, 66, -63, -57, -35, 39, -39, 47, -66, 50, 48, -36, 42, 67, 31, 22, -51, 26, -62, -60, 28, 50, 22, 34, -33, -17, 67, -25, 37, 0, 58, -9, -12, 70, 9, 27, 33, 43, -2, 41, 18, -32, -73, -18, -40, 33, -72, -16, -18, -61, -2, -66, 63, -56, 42, -46, 0, 31, 2, -39, -47, -16, 27, 17, -22, -42, -34, -67, -74, 37, 47, 17, -70, 49, 74, -37, 5, 75, 20, 62, -61, -58, 69, -74, -41, 33, -47, 34, -12, 28, 68, 17, -66, 19, -44, -15, 51, -5, -9, 52, -44, -37, -9, -41, -66, -11, -5, 14, -14, -60, 0, 0, -45, -6, -1, -10, -49, 25, -52, 13, -25, -59, -48, -16, 33, -19, 44, 8, 51, -40, -18, -71, -4, 46, -38, 5, -41, 32, -56, 21, 45, 19, -57, -75, -65, 16, -10, -40, -37, 11, 48, 14, 25, 73, 71, -17, -22, 38, 64, -47, 73, -31, -43, -9, -61, -8, 71, -28, -51, -63, 66, 67, 32, -67, 67, 40, 22, -21, 75, 61, 66, 45, -1, 15, 42, -8, 71, -56, -46, 58, -30, -51, -49, 1, 15, -37, 68, 9, 10, -61, 21, 0, -71, -25, 7, 71, -60, -47, -27, -63, -64, -37, 58, 8, 51, 22, -75, 47, 40, -46, 29, -68, -23, 53, 8, 67, -62, -1, 0, 24, 11, -54, -54, 15, -4, 26, 11, 9, 53, 57, 22, 64, -58, 2, -3, 68, -52, -3, 37, 61, 24, -12, 69, -75, -35, 1, 66, -23, 73, -10, -75, 9, 9, -56, -52, -72, 44, 32, 10, 21, 13, -44, 9, 30, 33, -72, 21, 55, -2, -18, 38, -53, 46, 31, -55, -67, -45, -65, -15, -48, -1, -17, 36, -70, 1, 58, -69, -31, 14, 17, 65, -50, 48, -4, 55, 4, 0, -2, -19, 71, 56, -57, -58, 26, 50, -39, 32, -71, -31, -60, -46, 43, -2, 64, 47, 74, 44, 53, -35, -18, -6, -48, 5, -35, 24, -15, 44, -54, 58, -51, -59, 36, -33, -43, -16, -61, -9, -59, -59, 35, -44, -31, 3, 27, -43, -26, 24, -75, -51, 64, -20, 19, -61, 61, 59, 38, -32, 25, 57, -52, 49, 71, 60, -62, -50, -34, -49, 16, -18, -33, -24, 11, 11, 52, -39, 41, -52, 60, 39, -28, 46, -56, 66, 60, -73, 47, 20, -30, -4, -1, -9, -33, -7, -25, -21, 18, 17, 5, -43, 72, 45, 8, 6, -19, -18, 42, -54, 5, 24, 61, 52, -8, -73, 41, -25, -71, 10, 68, -28, -71, -8, 38, -31, 58, -62, 23, 0, 28, -50, 32, 22, 71, -38, -48, -26, 19, 69, -7, -52, 15, -24, 74, -68, -22, 39, -18, -20, -29, -26, 27, -25, 39, -10, 20, 21, 1, -33, -54, -49, -9, 51, 48, -16, -64, -75, 33, 30, 67, -52, 52, 5, 0, 50, 12, 51, 11, 69, -44, 57, -35, 56, -43, -71, -32, 52, 25, 42, -59, 44, 68, 5, 18, 39, 64, 29, 37, 19, -19, 28, 43, -43, -43, -33, -69, 42, -60, 17, 33, -29, -1, 74, -50, 29, -73, -7, 3, 25, -42, 17, -8, -50, -53, -68, 64, -67, 34, 25, 28, -61, -24, -5, -28, 6, 37, -22, -29, 52, 69, -72, -54, -10, -74, -31, -57, -74, 35, 19, 25, 68, -40, -61, -59, -18, -54, -71, -11, 55, 28, -59, 69, -74, 11, -37, 5, -30, 17, 51, -56, 10, 53, -37, 73, 52, 7, -60, 54, -35, 32, 1, -43, 67, 13, -27, -28, 34, -24, 36, 11, -74, 52, 2, -75, -15, 39, 5, 30, -20, -21, 49, 63, -46, -65, 60, -70, 15, 73, 59, 55, 29, -18, -63, 20, 70, -17, 65, 26, 34, 25, -41, 33, -1, 35, 33, 59, -2, -39, 13, 51, 13, -15, 38, 42, -5, 20, 47, -66, 17, 29, 63, -32, -65, 75, 61, -72, -20, 51, 29, -63, -2, 62, 45, 73, 21, 3, 56, -57, 37, -8, 69, -26, 50, 29, -60, -33, -27, 60, -26, 63, 13, -39, -47, 22, -42, -62, 25, 14, 62, -24, 26, -15, -38, -5, -20, 56, 71, -42, 72, 32, 23, 65, -72, -3, 16, -59, 37, 62, -74, -64, 47, 14, -28, 75, -42, 4, -62, 56, -58, 73, -43, 43, -18, -8, -40, 35, -27, -46, 69, -33, 59, 14, -43, 63, -64, 46, -72, 46, 33, -73, 57, 4, 15, -48, 4, 48, 31, 15, 29, 48, 12, 59, 13, 68, -27, 46, 25, 19, 73, 16, 62, 57, -45, -59, 42, -36, 62, 43, -66, 17, 46, 67, -56, -15, -59, 21, -43, 47, -40, 59, 17, 45, 40, -48, 35, -62, 73, -15, 32, 71, 74, 16, 50, -47, 32, 16, -10, 17, -17, 0, -42, -47, -11, -25, 11, 5, 71, 44, -26, -47, 25, 66, 74, -10, -58, 31, 3, -63, -62, -43, -70, -63, 49, 55, -37, 3, -7, 29, -58, 50, -49, -24, -75, 15, 26, 12, -58, 20, -20, -9, 48, -73, -21, 46, -8, -4, 0, 70, 6, 13, -50, 12, 23, 72, -11, 62, -1, 56, 15, 17, 30, 41, 66, 30, -22, 14, -34, -7, -42, 19, 59, -69, 22, -38, 50, -64, 31, -26, -69, -41, 61, -46, 44, 8, -50, -44, -8, 22, -64, -69, -39, 41, 45, -51, -7, -55, 39, 33, 13, 70, -26, -6, 74, 69, 29, 47, -70, -18, -57, -66, 17, -72, -39, -17, 10, -14, 14, -74, -70, 25, -67, -33, -12, 51, -9, 55, 70, -48, 12, 7, -55, 59, 75, -57, 53, 28, 63, 56, -65, -69, 65, 25, -66, -52, -68, 19, 9, 22, 21, 14, -31, 27, 54, 31, 0, -32, 10, -6, -7, -54, 75, 13, -71, 74, 30, 55, 24, 17, 35, 32, 23, 22, -19, 31, 45, -13, -28, -24, -69, 68, 64, -27, 17, 42, -72, -60, -68, 13, 9, 1, 34, 6, -62, 37, 2, 41, 14, -49, -19, -28, 56, -72, 69, -40, 32, 37, 22, -71, -65, 26, 70, 74, 74, 12, 39, -73, 27, 46, 15, -42, -29, -28, 40, -17, -69, -36, -54, 20, -12, 2, 67, -31, 4, 59, 4, -40, 18, -52, -36, 28, 49, -43, 27, 45, 44, -12, 47, -7, -42, -15, 26, 3, 30, -12, 59, 36, 28, -71, -22, -60, 5, -30, -18, -67, -49, 61, -34, 44, -69, 4, -4, 53, 36, -55, 23, 4, 8, -8, 72, 40, 52, 20, -33, 6, -67, -52, -36, 36, -48, 18, 49, 32, 61, -44, 38, -64, -61, -71, 55, -54, 8, -27, 74, -34, -8, 21, 43, 75, -64, 39, 39, 63, -19, -72, -8, -11, -49, 29, -53, -23, -29, 70, -69, -46, -50, 45, -35, -38, 47, -58, -17, -23, -11, -20, 18, 56, 74, -15, 53, -66, -54, 15, 71, 2, 18, -13, 65, 43, -60, -64, -56, -15, -70, -52, 14, -47, 66, 53, -9, 37, 68, 47, -64, -19, -49, 27, -39, -50, -64, -61, -41, -45, 29, -48, 31, -31, 14, 20, -66, 28, 31, -49, -65, 35, -25, 24, 63, -35, -1, -24, -75, -8, -52, -64, 48, -28, 39, -68, -3, 48, -56, 30, -72, 46, 57, 34, -63, -6, -24, -53, -56, -71, -27, -46, 39, 21, 51, 25, 62, -25, -75, 60, 40, -54, 69, 12, -6, 32, 17, 64, 3, 36, 16, 4, 4, -4, -40, 17, 63, 11, 39, -69, 15, -66, -42, -21, 31, -67, -74, 15, -19, 75, -1, -55, -54, -10, 31, 13, -53, -28, -1, 23, -69, -62, -49, 10, 9, -14, -51, -6, 72, 63, 0, 9, 71, 31, 63, 26, 39, 62, -37, -57, 62, 35, -37, -70, -51, 67, 18, -31, -38, -61, 67, -32, -48, -58, 51, 34, 1, -75, -48, -5, 61, 25, -71, 56, -20, 65, 4, -58, 52, 42, -42, 38, 1, -6, 41, 26, -14, -19, 70, 23, -5, 60, 64, 21, 75, 37, -21, 1, 35, 5, 69, 21, -48, 73, -1, 6, 63, -72, 21, 37, 45, 54, -3, -29, -28, -38, 70, 33, 18, 64, -22, -65, 46, -36, 31, 46, -74, -67, -29, 34, 13, -38, -21, 38, -40, 54, -32, -55, 55, 64, 57, 24, 40, -22, 68, -63, 15, 62, 45, -45, 51, -54, -35, 21, -15, 72, -11, -16, -73, 33, -57, 15, 71, -5, -25, -45, -29, 17, -27, -50, 3, -46, 48, -32, 5, 40, -20, -56, 27, -53, -28, 0, -32, 12, -57, 27, 6, 8, -67, 8, -35, -49, -55, -40, 20, -4, -12, 64, -65, 36, -61, 13, 65, 62, 56, -8, 24, -42, 9, -25, -19, 56, 50, 22, -7, 67, -27, 72, -1, -20, 5, 37, 4, 25, 71, -52, -57, -17, -63, -47, -58, -51, 40, -71, -67, 20, -3, 32, 54, -70, -70, -43, 62, 55, 54, -23, 44, -50, -27, -33, 5, 51, -71, -67, -1, 75, -45, 15, -20, -35, 44, -3, -11, 8, 2, -5, -50, 74, -49, -74, -72, -44, -42, 63, -66, -63, -36, 53, -40, 11, -57, 38, -14, -55, 46, 58, -58, 74, -2, -3, -37, -34, 68, 25, 47, -6, -56, 70, -10, -31, 72, -9, -2, -46, -21, 7, -36, 16, -17, -1, -49, 1, -39, 11, 19, -70, -7, 36, -74, 66, -45, -37, -46, -55, 63, 74, 12, -70, 69, -74, -26, 65, -7, 47, -59, 45, -23, -21, -17, 33, 53, 10, -44, -63, -57, 50, -60, 11, 8, -61, 0, 36, -23, 27, 57, -37, 26, -7, -32, 17, -5, 15, 4, 61, -16, 20, 28, 34, 74, -65, -9, 50, 18, 22, 60, 36, -6, 75, -30, -74, -62, 43, 38, -11, -6, 17, 27, -58, -66, 70, 34, 2, 7, -38, -15, 66, 56, -63, 25, 54, -54, -62, 26, 39, 36, 10, -2, -46, 7, 41, -46, 19, 8, 65, -68, 75, 6, 32, -58, 15, 26, 51, -58, -45, -62, 0, -55, 69, 13, 43, 45, 32, 57, -6, -7, 15, -72, 66, 42, 9, 29, 71, -50, -39, 60, -45, -39, -10, 62, -24, -70, 10, -49, -55, 40, -38, 20, 58, -45, -45, 24, 74, 60, 5, -8, -22, -58, -7, -34, 59, 75, 71, 55, -51, -46, 39, -21, -12, -48, -37, 39, -45, 48, 66, -27, 10, -50, 66, -7, -19, -56, -59, -23, -72, 19, 44, -21, 36, -41, 21, 17, -41, 14, -4, -17, 43, -42, 36, -44, -17, 74, 68, 13, 45, 56, 61, -21, -69, 49, 45, -15, 68, 59, 37, 72, 2, 3, -25, -40, 37, 69, 53, 71, 7, -29, -23, -25, 2, -65, 4, 60, -69, -4, -5, 51, -23, -20, -45, -17, -48, 75, 43, -56, 59, 2, -60, -17, -71, -11, 17, 41, -18, -8, 35, 65, 36, -66, -38, -37, -56, 41, -53, -52, -41, 16, 75, 11, 69, -48, 67, -55, -51, 32, -35, -70, -42, -22, -11, -38, 42, -72, -74, -53, -7, 34, -64, -47, 43, -29, -9, 60, -64, 12, -68, -32, -50, -69, 53, -57, -44, 44, -36, -19, -1, 4, -14, 32, 57, 48, 68, 22, 51, 67, 44, -32, 25, 53, -5, -8, -52, 59, -26, -43, -7, -19, 0, 18, -14, -25, 37, 17, -56, -75, 73, 16, 2, -18, -28, -17, -46, -38, -73, -72, -47, 46, -31, 53, 21, 39, -33, 42, 23, 14, 74, -62, 71, -3, 32, -21, 47, -7, 69, 64, -9, 65, 4, 68, -29, 50, -27, 0, -66, -24, 3, -39, -56, 48, -64, 39, 9, -21, 5, -46, 66, 4, -32, 59, 74, 75, -38, 43, -10, -46, 30, 56, -57, -44, 48, -11, -72, -55, 62, -62, -6, -12, -26, 12, -42, -17, -25, 42, 35, 55, 72, 26, -19, -38, 9, -21, -39, 45, -55, 26, 74, 50, 6, -59, -72, -24, 3, -68, -6, -11, -57, 64, 52, -8, 0, -68, 48, 50, 50, 8, 27, 44, -42, -67, -70, 42, -15, -36, 9, 3, 65, 7, -23, -7, 21, -19, 42, -52, -14, -40, 11, 4, -52, -15, 69, 21, -7, 41, -7, -35, -27, -55, -67, 4, -49, -64, -31, 9, -25, 53, -63, -38, -15, -13, 28, -72, 41, -6, -48, -49, 29, 36, 30, 51, -55, 23, -6, 11, -13, 63, 51, 35, -70, 59, -36, -46, 70, 8, 38, -33, -17, 50, 4, 43, -38, -46, 45, -73, 23, 70, -46, -25, 30, 57, -50, 48, 3, 17, -16, 65, 4, -41, 22, 7, -59, 59, 36, -67, -9, -1, -24, 48, -29, 53, 13, 8, -68, -18, 9, 28, -24, 36, -73, -70, 15, -50, 54, -58, 43, -40, -69, -31, -6, 27, 52, 8, 10, 10, 17, 75, -69, 68, 47, -22, 43, -16, 59, 50, 42, -8, 3, -60, -50, 3, -54, 41, 29, 73, 58, -6, -45, 63, 36, 24, 14, 12, -43, -52, -55, 47, -55, -49, 39, 67, 2, 6, -24, -14, -21, -60, 51, 55, -45, -74, -18, -26, 42, -67, -31, 22, 0, -1, 9, -39, -54, -55, 46, -24, -33, 66, -53, -13, -60, 59, -21, 17, -13, 28, -75, 41, 41, 52, 18, 69, 53, -75, -34, 17, -69, 10, -37, 7, -68, 46, 43, -49, 64, 13, 2, -45, 2, 22, 16, 17, 3, 70, -42, 65, 20, -41, 29, -15, -67, -29, -24, 61, -31, 17, 0, -24, -48, 36, 56, -43, 4, 23, -17, -7, -42, 58, 21, 35, 2, -39, -24, -71, -47, 8, 69, 48, 40, 20, -45, 48, 65, 7, 31, -42, -54, -45, 7, -29, 64, -13, 3, -7, -66, 59, 59, -34, 41, 4, -75, -33, 41, -23, -31, 69, 58, -39, 40, 22, 56, 70, -6, 45, -1, -51, -74, 21, -23, 8, 67, -37, 71, -7, 31, -73, -24, 14, -32, -60, -59, -31, -20, 57, 19, 25, 48, 1, 61, 12, -53, 39, 7, 14, 7, -72, 36, 8, 22, -63, -60, 14, -27, -67, -71, -71, -64, -20, 16, -21, -7, 32, 21, 49, 11, -36, -4, -16, 38, -19, 71, 60, -58, 0, -4, 24, 4, -44, -46, -50, -34, -32, 37, 15, -24, 41, 17, -13, -56, -43, 40, 10, 63, -17, -17, -2, 21, 54, 55, -17, -43, 51, -32, -27, -27, 37, 70, 52, 69, -51, -75, -41, -8, 35, 49, 41, 1, -10, -47, 18, 21, 66, -48, 6, -29, 9, -74, 67, -15, 57, -25, 16, 30, 16, 64, -73, -23, 58, 53, -30, -71, 53, 3, -4, 12, -24, -38, -65, 40, -12, 26, -17, -24, 54, 64, 22, -15, 65, 12, 45, 46, 62, -15, 0, 0, -29, 1, 52, -48, -22, -55, -44, -45, 23, 26, 40, 74, 61, 49, 36, -29, -1, -57, 20, -25, -69, -34, 35, 72, 51, 3, 40, 37, 63, -37, -39, -43, 39, -64, -16, -61, -44, 15, -33, 54, -35, -69, 50, -52, 53, 9, -6, -23, 27, -62, 25, 32, -22, -15, 26, -47, 63, -10, 64, 48, 26, -53, -73, -13, -42, -14, 1, -13, -74, 43, -37, -36, 48, -64, -12, 25, 20, 55, -74, -29, 69, 27, -73, -29, -66, 28, -3, 70, -59, -15, 40, 42, 6, 43, -48, 39, -49, 28, -51, -48, -4, -13, -10, -32, -2, 51, 68, -60, 30, 68, -13, 21, 17, -13, 67, 24, -62, -13, 18, -46, 45, -20, 69, -25, -53, -55, -63, -26, 49, -39, -1, -33, 21, 62, 8, -58, 37, -2, -43, -10, -10, 19, -65, -71, -71, -75, 28, -58, -15, -32, -31, -46, 24, -38, 5, 44, -19, 17, -60, -48, 51, 13, -8, -4, -1, 75, 13, -41, -3, 44, 24, 61, -15, 32, 65, -11, 30, 16, 6, -61, 59, 48, -31, 5, -67, 49, -26, -11, -12, -13, 14, -37, 75, -70, 32, -1, -71, -32, 31, -1, -64, -21, -16, -4, -67, -28, 61, 39, 63, -11, 51, 44, -38, -56, -26, -30, 66, 21, 32, -24, -68, -32, 14, -68, -27, -31, 4, -25, 12, -41, 47, 21, 11, -44, -61, 17, 1, 75, -20, -14, -13, -46, -48, 22, -27, -1, 65, -38, -56, 19, 13, -50, 62, -50, -45, -43, -6, 34, 7, -72, 66, -24, 22, 1, 7, 36, -60, -70, 34, -4, -9, -55, 23, 19, 40, 71, -58, 29, -43, -40, -28, 46, -17, -44, 69, 13, -12, -13, -31, 68, -12, -41, -32, -66, 33, 49, 45, 48, 54, 3, -34, -32, 21, 64, 60, -15, 58, 75, -64, -63, -43, -19, 58, 15, 12, 51, -48, 73, -40, -6, 65, 21, 26, -42, 30, -17, -69, -2, -46, 58, 74, -7, -52, 20, -20, -68, -73, -38, -68, -63, -26, -36, -9, -45, 55, -74, -72, -71, 74, -38, -3, 64, 58, -53, -56, 13, 4, -52, -67, 33, -72, -69, -50, -48, 24, 5, -41, 25, 40, -36, 37, -61, 4, -50, -33, -19, -49, -30, -17, -50, 7, 55, -64, -12, -75, -45, 74, 4, -24, -69, -39, -21, -65, -16, 6, 35, 63, 39, -16, 27, -73, -57, 39, 4, -32, -70, 58, -5, -26, -34, 18, 54, -57, 29, -34, -57, 57, -36, 22, -43, -30, 56, 9, -21, -35, -62, -62, -50, 52, -5, 50, 52, 13, 14, -19, 54, 17, -37, -29, 64, 2, 64, 43, 19, 17, -67, 35, -4, -29, -18, 26, 14, -40, -40, 68, -2, -29, -72, 23, -55, -2, -2, 72, -67, -66, -25, 63, 26, 12, -42, 15, -62, -55, -20, 30, 35, -14, -10, -44, 32, 45, 57, -31, -71, -61, -39, 3, -15, -35, -50, 5, 36, 21, 0, 45, 30, 50, 30, -21, -14, 61, 67, -2, -70, -29, -48, 41, 30, 17, 72, -13, -14, 51, 29, -11, 66, 63, 67, -27, -50, -61, 52, 62, 36, -24, 29, -10, -52, -17, 42, 8, -32, 33, -70, -28, -72, -43, -65, 34, 48, -71, -57, -44, 55, 45, 20, 43, 32, 9, -61, 58, 22, 66, 42, -18, -36, -5, 45, -15, 51, 12, 68, -59, -31, 73, -12, -29, -47, -2, -73, 74, 2, -57, -48, -20, 63, 46, -53, 19, -21, -39, -1, -75, -51, -35, -20, -14, 33, -52, 47, 6, 33, 39, 23, 75, 35, -65, -30, 61, 7, -30, 59, -69, -12, -65, -14, -25, 54, 7, 68, -42, 41, -9, -44, 64, 30, 10, -26, -15, 33, -55, 67, -12, 58, 14, -13, 15, 22, 31, 0, -49, -75, -19, -42, -13, -11, 17, 37, -32, -52, 27, -1, 63, -59, 30, 51, 44, -38, -51, -47, 68, -32, -58, -20, -52, 29, 43, 38, -24, -2, -40, 2, -4, 16, 33, 58, -73, -25, 18, -30, -4, -31, 44, -17, -15, -3, -42, -47, 34, -19, -20, 27, 24, -3, -71, 45, -49, 47, 5, 0, -33, 40, 75, 39, -22, 33, 21, -20, -70, -39, 24, 1, 6, -10, 60, 64, 62, -60, -60, 19, -4, -5, -32, -58, 65, -28, 60, -60, -58, -11, 15, -16, -47, 13, -53, 4, -30, 42, 60, -27, -73, 6, 49, 6, 71, 31, -7, 56, 45, 8, -3, -35, -75, 38, -19, 65, -68, -35, -70, -51, 28, 18, 7, 54, -45, 27, -17, -2, -7, -35, 46, -6, 46, 18, 73, 39, -27, -10, 19, -58, 71, -60, -19, 71, 51, 35, 61, 59, 73, 64, -68, 25, 4, 14, 4, 33, -34, 60, -45, 32, -51, 75, -52, 68, 17, -54, 31, 63, 9, -27, -72, 3, -14, -16, -2, -38, -59, -19, -55, -62, -33, -48, 37, 47, 40, -37, 2, -70, -53, 30, 35, -31, 29, 59, -39, -32, -73, 65, -46, 9, -38, -43, -64, 22, 14, 8, 59, 30, 64, -72, 41, -46, -47, 2, 74, 68, 38, 0, 71, 60, -48, 29, -49, 57, 12, -13, -53, 12, -25, -24, -55, 12, 6, -45, -42, -56, 38, -61, 47, 24, -58, 13, 53, -31, -63, 51, -39, 49, -27, -45, 33, 1, 59, 60, -20, -7, -31, 0, -71, 19, 50, -53, -46, -20, -23, -15, -2, -61, 0, -31, 39, 15, 55, 14, 59, 66, -12, -57, 39, 36, -27, -6, -41, -46, -24, 14, 20, 19, -63, 24, -38, 62, 44, -11, -34, -54, 50, 39, -42, -28, -69, 70, 62, 59, 9, 44, 49, 70, 62, 10, 28, -43, -71, 63, -14, -22, -1, -70, 72, 11, 27, -43, -3, -5, 19, 37, 14, -9, -2, 48, 38, 4, 40, 23, -12, -27, -9, -41, -35, -23, 45, 69, 9, 47, 56, 68, -53, -21, 71, -58, 66, 22, -26, -15, -61, 68, -54, 27, -16, 20, -1, -56, -54, -37, 42, 7, 10, -45, 42, 50, 7, 9, 43, -62, -22, 21, -70, -2, -75, -75, 15, 64, 20, 62, -27, 33, 53, -7, -16, -39, -65, 56, -22, -44, -59, -57, 39, 26, -27, 3, -1, 56, -66, -36, 67, -15, 61, 71, 58, 59, 69, -4, 45, 14, -18, -60, -31, -41, 8, 26, -7, 18, 6, 47, 50, 22, 63, 11, -29, -40, -64, 43, -62, -57, -69, -70, 3, 65, -75, -17, 46, 69, 54, 15, 5, -41, 31, 47, -7, -37, -3, 62, 55, -73, 31, 27, 23, 18, -38, 67, 51, -29, 34, 65, -11, 38, 68, 67, 28, 66, -28, -2, 57, -51, -62, -15, -17, 42, -44, 51, -71, 27, 35, 59, 29, -12, 10, -26, -72, 45, -35, 55, -60, 74, 42, 4, 37, 32, -7, -13, 20, 39, 58, 1, 63, 69, 59, -32, 35, -62, -57, 38, 40, 52, 21, -9, -38, -46, 41, -34, 72, -72, -55, -63, -73, 60, 14, 37, 14, -70, -54, -42, 42, -72, 34, 27, 71, 16, 70, 30, 29, -65, -8, -7, 62, -64, 59, -51, -37, 22, -12, -41, 26, 6, -31, 26, -10, 57, -13, -72, 60, 6, -41, 26, 7, 68, -23, 2, 6, -29, -45, -41, -19, 20, 27, -34, 31, 9, -12, 69, -45, 51, -49, 56, -21, -5, 6, 44, -24, 66, 45, -40, -6, -72, 59, -74, 69, -40, 1, 0, 4, 31, 34, 59, -24, -16, -51, -71, 66, 10, 72, -55, -17, -53, 75, 37, 15, 3, 3, 65, -6, -28, -53, 63, -27, -69, 62, -36, -36, -12, 37, 44, -59, -6, 27, -8, 53, 49, -5, 43, -19, -9, 61, 39, 11, 60, 0, -50, -12, -73, -61, 55, -28, -40, 40, 18, -34, 27, 57, 3, -61, 19, -29, -47, -63, 71, 21, 63, 42, -60, 30, -53, 4, 13, 61, -61, -2, -15, -36, 59, -15, -23, 36, 30, 12, 0, -28, 51, -49, -46, -22, -37, 48, 23, -8, 58, 16, -65, 45, -17, -52, -3, 5, 27, -66, -11, 41, 5, 47, -71, -14, -43, -21, -54, 62, 64, 22, -43, 37, 46, -14, -60, -68, -44, 36, -1, -64, -24, 7, 56, 32, 30, -23, -40, -19, -16, 24, -54, 63, -5, -52, -27, 25, 1, -5, 10, -11, -61, 42, -49, 60, -50, -36, 65, -19, 73, -14, -8, -27, 68, -30, -72, 20, 20, -37, -75, -74, 62, -56, 64, -21, -34, -40, -73, 42, 28, 12, -47, 42, -24, -21, 24, 1, 16, 14, 55, 13, 75, -31, 60, 68, 14, 63, 10, -44, -52, 11, -43, -68, 28, -54, -14, 69, -21, -12, 33, -69, 73, 62, 48, -27, -37, -4, 47, 55, -68, 26, -10, -68, 68, -26, 73, 6, -41, 7, 35, -18, -60, 68, -11, 42, -64, 49, 35, -10, -41, -9, -4, -43, -23, -34, 3, 13, 35, -27, -10, 43, 72, 56, 48, 65, -46, 43, -7, -13, -28, -47, 44, -14, -57, -44, -48, -46, -71, 60, 17, -37, -25, -63, -7, 25, -24, 72, -37, -65, -33, 26, 53, -37, 6, 23, -48, 34, -10, 19, -55, 36, 47, 62, -54, 65, -58, -27, -59, -54, -43, 31, -15, 6, 43, 51, -45, -59, 45, -9, -49, -64, -60, -73, -25, 21, 25, 0, -23, -62, -57, -5, 47, 63, -18, 68, 50, -1, -37, 66, 19, -5, 21, -74, 74, -14, 52, -48, 2, 22, 16, 27, 33, 31, 29, -70, -23, -24, 6, 27, -13, 22, -53, -42, 10, 4, -50, -16, -75, -12, -27, 19, 57, 67, 20, 53, -22, -3, -71, 53, -57, 21, 4, 49, -24, -45, 53, 26, 5, -19, -22, 67, -73, 0, -52, 10, -74, -29, 70, -74, 35, -35, 21, 14, -44, -35, -9, 7, 35, -6, -15, 51, -61, 62, 25, -12, -60, 0, -61, 20, 56, -10, 9, 56, 63, 32, -9, 64, -72, -17, 65, 36, 23, 10, -28, 54, 49, 36, -14, 8, -46, 44, -16, -34, 28, -69, 30, 43, 4, 42, -15, -16, -44, 70, -36, -57, 24, 30, -71, 25, -65, 69, -15, 33, 2, 30, 10, -25, -9, 69, 56, 18, 35, -38, 60, -13, -34, 12, -45, 45, -22, 13, -47, 7, 7, -9, 23, -46, -57, 27, 54, -46, 20, -38, 62, -56, 67, -6, -6, -20, -13, -27, 74, -54, 10, 56, 9, 52, -8, 37, 21, 45, -26, 48, -26, 55, -37, 72, -67, -21, 23, 60, 8, -35, -54, -5, -15, -64, 64, 52, -9, -26, -51, -13, -5, 33, -35, -74, 9, 32, 36, -48, -1, -65, 73, 48, 63, -42, 42, 71, 13, -13, 55, -55, 28, 75, 13, -65, -65, 0, 60, -1, 49, -66, 60, -34, 40, -51, -34, -27, 55, -74, -2, -22, -66, -4, -51, 72, 27, 66, 65, -36, -22, 43, -17, -72, 40, 71, -64, 48, -7, 71, -29, -34, -73, -47, 6, 42, -24, 45, -63, -45, 44, 11, 8, 54, -71, 32, 48, 31, 21, 36, 69, 74, 1, -26, 75, -35, -31, -65, -63, 36, -70, -19, 75, -67, 10, 5, 50, 61, -28, 63, -62, -59, -4, 21, 68, 0, -24, 38, -47, 72, -4, -56, 68, 72, -7, 67, -39, 36, -74, -29, -4, -69, 28, -5, -61, -40, 74, 63, -57, -30, 48, -44, -16, -32, 50, -24, 41, -50, -63, 69, -56, 8, -64, -64, 5, 4, -73, 39, -38, -72, -65, 31, -67, 36, -49, -55, 71, -53, -68, -64, -10, 55, -33, 50, -55, -59, -52, 61, -35, -40, 55, -16, 44, 64, -4, -29, -10, -4, -66, 28, -2, -58, -17, 6, 53, 7, 24, 46, 27, 30, 57, -58, 7, -54, 65, 28, -39, -63, 13, 1, -29, -10, 58, -63, -22, -24, -17, 44, 48, -10, -6, -30, 6, 52, 49, -17, -18, -3, -48, -67, -49, -69, -50, 34, -47, -61, -14, -13, -50, 72, 63, -4, -13, 43, 6, 38, -56, 64, 4, 67, -24, 73, -41, 57, 48, -68, -37, -46, 2, -10, -38, 29, -6, -14, -15, 20, -2, 44, -69, 21, 40, 67, -61, -51, 35, 20, 61, 54, 8, -11, 45, 58, -13, -74, 39, -41, -67, -74, -14, 8, -11, 23, -41, 57, -69, 19, 1, 5, -15, 6, -52, -52, -3, -37, -30, -44, 58, -45, -68, -11, 20, 52, -29, -71, 51, -68, -37, 59, -68, 24, -8, -6, -31, 26, -25, -26, -32, 50, 52, 26, -20, 75, 49, 52, -38, -56, -69, -55, -26, -62, 9, 67, 64, 53, 71, 39, 60, -44, 21, 65, 55, -63, -16, -53, 36, 34, -4, -74, 8, -28, 28, 63, -29, 1, 38, 7, 18, 44, 27, 68, 57, -42, 59, 45, -65, 53, 7, 68, -67, -48, 58, 62, -36, -34, -67, 73, 73, 2, 73, 4, 47, 23, -9, -60, -54, -49, 22, 40, 70, -27, 30, 50, 4, 11, 19, 12, -12, -52, 5, -3, -25, -15, -17, 12, 26, -11, 10, 21, 66, 5, -51, 35, -48, 14, 50, -27, 40, -3, -65, 33, 43, 40, 7, -28, -26, -52, 59, 37, -28, -14, -42, 22, 46, 14, -41, -6, -73, 42, -62, 66, -31, -38, 25, -4, 49, 0, 42, 12, 70, 53, -31, 37, 15, 49, -69, 64, 72, 64, 24, -34, -26, 55, 64, -57, -6, -55, 10, -6, 60, 23, -15, -47, 61, -66, 24, 32, 7, -12, -32, 1, -37, 12, -39, 52, -15, -33, 40, -20, -45, -14, 21, 3, -34, 7, 21, 35, 25, -45, -47, 9, 54, 11, 37, 37, 19, -17, -7, -50, 45, 37, 25, -68, -29, 61, 59, 30, -48, 22, -66, -19, -68, 28, 57, -27, -40, 2, -70, 60, 30, -43, -8, 6, 43, -47, -35, -14, 12, 32, 10, -19, -7, -41, -14, 37, -56, -32, -9, -31, 65, -2, 23, 70, -49, 4, -34, -16, -72, -29, -34, 32, 3, 33, -38, -31, 62, 1, 30, -4, -43, -36, 50, 23, -4, -42, -16, 13, 1, 49, 58, -12, -29, 3, -17, -5, -68, 24, 52, -67, 68, -57, 40, -6, 51, -73, 38, 35, 1, -10, -47, 33, 30, -73, -20, -52, -41, 37, 37, 35, 10, 17, -52, 55, -56, 4, -28, -51, -50, -51, -42, -60, -33, 73, 9, -60, 73, -29, 51, -2, 37, -72, -47, -11, -71, 6, 10, -37, -32, -29, 71, 51, 61, -59, 28, -72, 20, -75, -48, 43, -51, -17, 59, -9, -21, -8, 4, -24, 37, -21, 48, -4, -19, 74, 58, -15, 5, -8, 21, 48, 39, 16, 23, 22, 33, -26, 25, -25, -26, 51, -57, -2, -42, -74, 62, 12, -9, -10, 62, -50, 43, 32, 21, -52, 30, 3, 8, -41, 71, -47, -71, 32, 42, 26, -22, -1, 75, -74, 50, -27, 52, 68, 44, -66, 67, 30, 20, -20, -58, 6, 4, 60, -38, -53, -68, 65, 26, 13, -51, 19, 39, -47, -27, 6, 52, 24, -71, 51, 25, 54, -52, -1, 44, 67, 9, 33, 19, -49, -64, 37, 32, 15, 19, 67, 37, 27, 54, -15, -38, -75, -74, -74, -48, -28, 7, -72, 70, 9, 55, 17, -14, -75, -59, -46, 66, 23, 61, 9, 49, 72, -32, 3, 9, 63, -8, -32, 12, -30, 27, 49, -29, 28, 48, -2, 74, -21, 1, 68, 64, -22, 9, -26, -21, 23, 1, -31, -30, -14, 51, -59, -20, -56, 19, 62, -71, -67, -45, 14, -21, 57, -15, 23, 7, -42, -57, 5, 12, 17, -5, -2, 71, -71, 45, -28, 27, -29, 14, 71, 30, -11, -64, -67, 6, 31, 70, 10, 37, -53, -52, -62, -72, 9, 36, 11, 40, 52, -62, -24, -6, 9, 48, -13, 11, 17, 34, -38, 61, -28, -45, 16, 34, -33, 22, -35, 71, 16, 48, 32, 37, 72, 46, 40, 3, 4, -27, -33, -19, -15, 16, 48, 69, -12, -41, 4, -72, 66, 39, 64, -40, 70, 2, 69, -41, -52, -44, -48, 38, -71, 59, -1, -75, 27, -39, 1, -44, 8, 41, 10, 68, -19, -18, 59, 43, 14, -13, 44, 4, -52, 30, 37, -60, -43, 30, -26, -22, 60, -1, -62, 64, -17, 10, 62, -68, 45, -13, -39, -23, -50, 46, -31, 4, -50, -48, -29, 39, 12, -63, -35, 33, 43, 75, 49, 73, 28, -55, -27, 12, 20, -15, 0, -75, 70, -14, -68, 39, 46, -31, -62, 71, -63, -20, -1, -37, 5, 44, 75, -59, 56, -37, 48, 21, -40, 21, 16, 63, 39, 65, -1, -19, -28, 74, -19, -34, -18, -13, -72, -48, 31, -61, -53, 41, -5, 20, -72, 75, -12, -74, -61, -34, -38, 62, 61, -3, 5, 1, -15, -32, -12, 57, 25, 35, 56, -72, 75, -40, -10, -75, -12, -55, -61, 8, 62, 9, -48, 63, 7, 13, 62, 19, 55, -54, 5, 40, 19, -66, -37, -74, -25, 27, 58, 73, -16, 36, -74, -17, 70, -9, -17, -18, 10, -4, 63, -6, -73, -62, -21, 9, 26, -34, -50, 3, -15, 30, -35, -74, 37, 4, -73, -65, -47, 59, -68, 12, 17, -67, 69, 9, -2, -24, 66, -68, 45, 52, 1, 48, 65, 55, -21, 13, -57, 5, -61, 4, -43, -21, 5, 70, 56, 6, -73, -67, -13, -66, 19, -74, -59, 12, 11, 14, 61, -1, 21, 31, -27, -56, 3, -38, 74, 55, 49, -60, -16, 63, 17, 17, -36, -54, 9, -55, 25, 11, -49, -66, 18, 45, -66, 34, -21, 20, -28, -35, -59, 66, 69, -10, -66, -6, 25, -69, -27, -4, -54, 31, -17, 36, -30, 21, 55, 54, 39, 5, -13, 65, 12, -73, 33, 21, 37, -66, -37, -69, -26, -20, 73, -33, 43, -71, 34, -10, -67, -68, 62, -48, 38, -33, 63, -70, 63, 43, 57, 26, -30, -32, 14, 57, -30, -29, 1, -71, -20, 39, -64, 28, -59, -69, 68, 59, -65, 27, -28, -56, 32, -42, -29, -6, 0, -41, -3, -12, -74, -22, -64, -31, 21, 25, -50, 64, 69, 26, 67, -26, -12, -73, 75, 4, -67, 67, -14, -59, 16, 33, -42, -28, 66, 5, 39, -12, 37, -40, 49, 36, 13, 61, -71, -44, 10, -48, -57, 2, 54, -66, 51, -34, -66, 48, 43, -60, 37, -49, -44, -22, 59, -12, 23, 47, 66, -13, -42, 27, 22, -69, -15, -42, 67, -13, -11, 0, 14, 5, -74, -10, 14, 50, 29, 23, 20, -3, 36, -19, 23, 68, 32, 5, -20, -20, -26, -32, 42, 7, 70, -14, 14, -23, 19, 3, 39, -69, -75, -25, 11, -74, 41, -52, 49, -8, 44, -7, 62, 5, 48, 8, -5, 4, -63, 48, 59, -16, -60, 25, 67, -68, -64, 3, -16, 28, -70, -55, 34, -69, -5, -32, -70, -42, -11, 55, 26, -43, -30, 10, 35, -58, -58, -46, 22, -46, 75, 5, 12, -61, -47, 3, -54, -38, -70, 3, 65, -67, 21, 22, -61, -61, 65, -57, -28, -24, 73, 71, 8, -35, 6, -34, -19, 23, -5, -73, 51, -7, 5, -13, 7, 31, 63, 27, 68, 68, -48, 56, 74, 49, 2, -62, 63, -11, -44, -43, 40, -49, -47, -30, -11, 32, 11, 45, -23, -71, 45, -50, -3, -27, 12, -74, -72, -3, 28, 70, -11, 54, 50, -14, 27, -26, -1, 12, 38, 28, 44, 0, 52, 70, 43, -37, 24, -21, -67, -74, -19, 51, -49, 53, -52, 37, 54, -50, -42, 5, -56, 21, -17, 69, -69, -68, -35, 3, 19, -75, -47, -13, 0, -71, -20, -35, -35, -72, 17, -29, -73, 73, -53, -46, 50, -30, 64, 27, -5, -54, -44, 12, 42, 12, 5, 46, 19, 43, -27, -38, 43, 1, 22, -35, 3, -74, 6, 44, -72, -53, -61, -70, -55, -41, -43, 68, 5, -55, 17, 73, -33, 46, 10, -69, -18, -63, 53, 74, 56, -52, -40, 21, 23, 56, 62, -50, 57, -8, 67, 58, 14, -71, 64, 32, -37, -55, 23, 41, -34, -36, 37, 6, -67, -31, 10, -10, -21, -13, -11, -43, 9, 22, 54, -44, 2, 40, -21, -18, -44, -31, -38, 43, -27, -50, -2, 9, -31, -55, -27, 8, -18, -66, -62, -10, -24, 21, 56, 30, -67, -33, 63, 15, 62, 41, 46, -13, 5, -53, 42, 34, -9, -72, 1, 37, -48, 74, -29, -4, -59, 19, -74, -1, 26, -63, 64, -74, 33, 42, 29, 39, -67, 16, -22, 69, -21, -54, -20, 59, -31, -54, 15, 35, -53, -59, -3, -26, -63, 41, 43, -46, -18, 44, 28, -68, 54, 14, -69, 12, -19, 35, -25, -13, -26, 27, -20, 28, 48, 35, 10, -59, 54, -51, 50, -74, -35, -31, -27, -24, -66, -59, 3, -9, 58, -47, -4, 35, 42, 2, -29, -53, -41, 19, 10, 8, -30, 65, -41, -59, 23, 44, -45, -1, 68, -71, -2, -44, -27, 47, 5, -20, 61, -68, 46, 41, -40, -34, 0, 75, 41, 44, -55, -75, -12, 30, 6, 31, 17, 38, 47, -38, 6, -75, 37, -1, -71, -43, 28, -24, -72, -43, 31, 62, -38, 0, 26, -3, 41, -50, -6, 5, 70, 14, 3, -20, -32, -67, -65, 59, 47, 56, -57, -25, 56, 55, 47, 58, -63, -1, -42, -62, 29, 63, 74, 66, -13, 24, -15, -50, 47, 55, 30, 41, -9, -43, -57, 33, -36, -46, 16, -67, -68, 34, -17, 63, 12, -47, 43, 22, 25, 75, 33, -21, 62, 31, -33, -29, -23, 28, -6, -51, 5, -51, 63, 69, -21, -69, 26, 18, -42, -36, 24, -35, 72, -70, -50, 8, -42, 68, -48, 58, 67, 58, -39, 51, 14, 2, -56, 66, -48, 14, -63, 30, 38, -75, 23, -61, -69, -26, 31, -36, 13, -21, 4, 7, -16, 27, -63, 15, 19, -36, -2, 9, -53, 32, -16, 34, -42, 4, 22, -15, -60, 35, -63, 53, 33, 36, 65, 39, -68, 20, -73, 18, 73, 4, -50, -21, -45, -38, 70, 47, 0, -10, -20, 20, -54, 38, -22, -22, -34, 73, 36, -19, 30, 49, -44, -13, 7, -57, -50, 14, 39, -50, -44, 34, 27, -19, -63, 57, 17, -69, 27, -59, -6, -69, 36, 16, 44, -64, 69, -68, -69, 27, -14, 37, 0, 15, -54, -69, 34, -30, 18, -5, -5, 50, -47, -55, -47, -37, 75, 43, -32, 26, 59, 37, 31, 17, -25, -1, 26, -34, 5, 33, 69, 66, -8, -9, 4, 13, -4, -38, 58, -62, 30, -24, 61, 56, -6, -61, -57, -7, 57, -14, -56, 39, -54, 50, -22, -4, -29, -71, 38, 51, 35, 31, 40, -49, -54, -32, 37, 17, 3, 20, 31, -43, 69, 14, -63, -13, 28, -45, 53, 8, 15, 72, -31, 36, 44, 20, -44, -62, 22, 69, 62, -19, 22, 26, 5, 42, 69, -33, -17, -6, 60, -64, 26, 51, 26, 38, -38, -24, 67, -61, 57, 4, -66, -52, -36, 51, 44, -7, 64, -10, -15, 51, 47, -69, -1, -26, 46, -9, 16, -48, 60, 0, -39, 11, -25, 60, -29, 10, -39, -40, 23, -60, 39, 30, -36, -73, 5, -68, -6, -8, -5, 54, -35, -36, 58, 39, 14, 29, -48, -46, 56, -63, 28, -61, 21, -75, 75, 65, 9, -40, -50, -44, -27, 64, 61, 12, 65, -12, 17, -17, 55, -65, -41, -58, -26, -61, 55, 63, 43, -69, -60, 21, -59, 41, 36, 35, 39, 35, 25, -28, 68, 50, 1, -35, 36, -16, 51, 25, 48, -10, -70, 25, 0, -36, 41, 48, -21, 20, 33, -56, 24, 48, 39, 41, 11, -3, -2, -25, -46, -53, 20, -54, 70, -56, -16, 31, 3, -43, -22, -27, 21, -16, 74, -57, 23, 39, 66, 75, -19, 24, -56, -71, -6, 56, 43, -72, -23, -34, -24, 6, -14, 71, 25, -19, -61, -69, -66, 16, -38, -13, 64, 58, 46, 62, -75, -8, 23, 65, -9, -74, 11, 8, -69, -71, -14, 47, -70, 38, -65, -19, -34, -5, -25, 66, 51, -11, 71, 58, -71, -43, -31, 69, -61, -60, 53, -63, 5, -1, 75, 69, 0, 10, 2, 4, 13, 63, -26, 18, 24, -16, 75, 65, 52, -26, 54, 25, 36, 47, 7, 39, -72, 52, 30, -60, 65, 7, -50, -6, -72, -50, -13, 4, 35, 62, -68, -30, 48, -21, 64, -4, 39, 61, -17, 13, -43, -41, -37, 68, -70, 45, 29, -67, 19, -17, -54, 8, 64, -28, 75, 67, -5, -15, -7, -46, -31, 1, 0, -61, 55, -14, 10, 16, -29, 67, -46, 3, -50, -10, -7, -44, -41, -53, -38, 52, 3, -18, -18, -9, 27, -18, -19, -54, 40, 49, -27, -69, -28, 46, -54, -50, -44, 29, 39, 0, 20, 66, -75, 44, -20, -8, 73, 13, 14, -43, -11, -61, 14, 46, 4, -35, -50, 60, -16, 63, 33, 33, 70, -72, 3, -62, -47, 33, 42, 67, -43, -15, 58, -44, -47, -40, 23, -52, 48, -41, -20, -39, -27, 68, -70, 52, -45, -45, 36, 15, -57, -8, -28, -65, -5, 48, -52, 23, 3, 63, 12, 34, -28, -8, 65, -2, 28, 12, 21, 0, 46, 75, 35, -59, 65, 40, 69, -56, 68, 27, 34, -65, -57, -72, -55, 11, 50, -34, -44, -23, -46, 44, -65, -1, -40, 73, 73, 61, 9, 16, -16, -23, 13, -57, -6, 2, 56, -13, 22, 48, -64, -22, 57, -47, -20, 75, 39, -48, -34, 71, 2, -7, 39, 11, 67, 72, 8, 62, 58, -58, 3, -34, -8, -62, -18, 61, 16, -38, -30, -40, -68, -18, 11, 62, 10, 64, 62, -29, -60, -50, -34, 16, 18, -73, -49, 9, 75, 34, -6, 55, 49, 70, -55, -34, -68, 2, -49, 21, 37, -5, 56, 42, 50, -10, 29, -18, -24, 15, 28, -10, 40, 70, -70, -18, 70, -44, 64, 69, 63, -20, 48, 37, -26, 66, -75, -18, -8, -51, -75, -49, 19, 57, 69, -7, -31, 22, 50, 20, -41, 1, -66, 74, -5, -61, -22, -13, -32, -36, -19, -46, 20, -49, 66, 69, -60, 64, -27, 7, -63, -26, 32, 30, -47, 25, -55, -5, -31, 69, -61, 3, -6, -53, -1, 62, -41, 52, -27, 1, -62, 27, 30, 33, 52, 18, 25, 67, 6, 71, -4, 16, -33, -48, -30, -7, 50, -9, 63, -57, -18, -75, 19, 51, -53, -58, 37, -21, 67, -68, 55, -70, 35, 9, 36, 9, -51, -15, 0, 30, -21, 71, -29, 21, -54, 14, -61, 71, -73, 75, -63, -16, 75, 29, -41, -54, 47, 69, -1, 36, -74, -22, 41, 34, 61, 2, -33, -66, 60, 40, 38, -37, 35, -69, 58, 56, 20, 72, 50, 23, 69, 60, -71, 69, 13, -38, -63, -18, -45, 11, -57, -46, 63, 57, 61, 48, -17, -50, 55, -32, 65, 17, 4, 23, 23, -14, 1, -32, -20, -27, 64, -26, -43, 66, -33, 44, -48, -23, -50, -19, 64, -34, 8, 51, -52, -8, 21, 4, 17, 0, 45, 5, -58, -26, -48, 38, 33, 26, -72, -62, 75, 67, -15, -44, 58, 25, 73, -68, -74, -54, -12, 65, -13, 70, 38, 8, -14, -19, -63, -73, 57, 57, 5, 72, -47, 32, 34, 62, -19, 38, 73, -20, 27, -18, 11, 7, -69, 9, 15, -68, 28, -75, 71, -61, 70, 31, 21, -22, -63, 33, -21, 67, 12, 59, 63, 41, 14, 19, 27, 70, -21, 24, -26, -69, -72, 58, 11, -66, -11, -50, -61, -59, -51, -68, -44, -59, 39, 50, -5, 49, 7, 49, 40, -59, 32, 25, 57, -30, -32, 6, -38, 23, -48, 11, 27, -45, -6, -38, -38, 56, -14, -23, 73, 10, -16, -49, 24, -55, -75, -57, 69, 5, 67, 33, 21, 22, -20, 3, 67, 24, -69, -46, -31, -41, 38, 71, -11, -46, -45, 25, -65, 14, -74, -68, -54, -17, -42, 46, 4, -44, 64, -5, 36, 54, -49, -19, 0, 6, 57, -11, -46, 64, 18, -4, -53, -21, -11, 9, 8, 20, -42, 18, -42, -43, 23, -20, 16, 56, -52, -58, -66, -64, 10, 45, 65, 36, -51, -13, -33, -70, 52, -6, 69, -8, 66, -62, 46, -23, 23, -21, 72, 54, 70, -47, -64, 18, 6, 25, -4, 29, 40, 6, 38, -26, -27, 26, -65, -3, -63, -25, 3, 64, 44, -6, -19, 32, 8, -51, -66, -45, 3, -72, -67, -4, -46, -58, -62, 33, 42, 9, -16, 4, -63, -53, 54, -14, 46, 62, 58, 58, -39, -17, 47, -73, 53, -50, 33, -15, -26, 40, 13, 51, 43, 19, -29, 71, 37, -16, 28, 1, 66, -63, -70, -72, -43, 57, -13, -73, 43, -31, 60, -72, 26, 29, -72, 1, 52, 36, 61, -49, 0, -4, 75, -34, -61, -30, -39, 49, 27, 62, -27, 15, 72, -22, 18, -47, -43, -71, -45, 75, -28, -62, -75, 71, 40, -72, -4, 17, 38, -21, 41, -38, 50, 40, 1, 62, -68, 35, 36, 32, 22, -67, -29, 18, -16, 63, 47, 16, 67, 75, 15, -39, -65, 13, -44, 51, 16, 25, -8, -24, -72, -45, 14, 53, 68, -63, 40, 75, 48, -2, 29, -6, 4, 75, -66, 63, 62, 54, 3, 52, 54, -60, -65, 64, 28, -33, 37, -34, 67, -47, 18, 69, -19, -46, 46, -27, -34, 8, -30, -64, -72, 74, 3, 7, 72, 13, -6, 56, -9, 70, 32, -33, -68, 41, -46, 33, -68, 66, 75, 72, -58, 15, 65, -4, 42, 34, 45, -70, -36, -61, -58, -32, -64, 20, 48, -68, -43, -33, 63, 22, -41, 18, 62, -33, -17, -62, 75, -12, -71, 72, -18, -56, 9, -28, 15, -25, -72, -18, -19, -35, -3, -2, 8, 6, -60, -19, 13, -29, 21, -2, 68, 55, -62, 52, -56, -6, 66, -58, 57, 68, -62, -38, -66, 23, 7, 24, 71, 10, -71, -26, 50, -1, 47, -19, -71, 61, 35, 15, -44, -20, -65, -54, -43, -51, 73, -25, 18, 61, -8, -2, 53, 5, 33, 62, -50, -36, 9, -56, 47, 13, -7, 21, -64, -37, 75, -60, -52, 34, 28, -23, -64, 38, -2, -33, 62, -7, 17, 3, -23, -67, 74, -46, 11, 31, -61, 35, 68, 23, 54, 39, -42, -31, -18, -33, 7, -18, -20, 28, -62, -68, -71, -52, 45, 0, -10, 30, 67, -69, -45, -32, -63, -47, -3, 23, 57, 9, -20, 47, -46, -42, 10, -13, 3, 67, 29, -68, -29, -67, 36, -17, -62, 40, 6, 59, -37, 69, 13, -46, 73, 41, -3, -66, 69, 67, 30, 48, -1, -65, 19, 28, -34, -49, -60, 44, -60, 42, 50, -13, 49, 10, 43, 62, -28, -29, 45, 10, -36, -20, 37, -39, -55, -44, -30, -64, -54, 75, 57, 20, -68, -2, -28, -26, 24, -15, -58, 38, -48, 65, -53, 74, -1, 65, 60, 45, -40, 30, -23, -1, -68, -61, 33, -49, -32, -73, -40, -11, 75, -58, -69, -68, 13, -23, -19, -40, 35, -4, 73, 60, -14, -56, 58, 58, -69, 43, 27, -36, -5, -71, 36, 2, -59, -7, 26, -16, -7, 62, 47, -8, -74, 51, -3, 12, -48, 51, 47, 63, -28, 42, 47, 31, 59, 30, 13, 65, -5, -37, -47, 65, -33, 64, -11, -19, -21, -60, 40, 47, 75, 9, -38, 74, -15, 34, 10, 10, 10, -20, -3, 55, -54, -33, 8, -70, 70, -57, 68, -11, -19, -56, -22, 21, -70, 40, -74, -15, 53, 40, -46, 52, -27, -9, 48, 31, -50, -17, -34, 33, 36, 38, 10, 57, -73, -58, 60, 72, -40, 51, -17, 17, 68, 34, -40, 73, -1, -38, -20, -24, -74, 10, -49, -28, -75, 72, -72, -52, -21, -31, 54, -63, -71, -12, 68, -68, 3, 52, -74, 37, 25, -15, -24, 17, -59, 11, 13, 15, 48, 66, 65, 47, 0, -62, -56, -1, -66, -53, 20, -13, -9, -1, -1, -7, 60, -9, 0, -12, -34, 0, -51, 64, 58, 0, 4, 74, -65, -59, 12, 57, -69, -1, 28, 5, 12, 47, -72, 19, 67, 21, -70, -20, -56, 3, 49, -71, 67, -29, -8, -43, 46, 14, -56, 26, -62, 23, 25, -54, 39, -41, -73, 43, 33, 31, -30, -31, 0, -29, 63, -8, 68, 67, 45, -64, -6, 18, -62, -15, 63, 3, 16, 31, -59, 35, -18, -48, -20, -71, -26, -57, -37, -24, 59, 71, -71, -46, -36, 3, -2, -51, 68, -10, -62, 37, 0, 5, -22, 13, 64, -35, -59, 4, 71, -43, -39, -25, -15, 16, -21, 32, 32, 17, -70, 13, 12, -65, 42, 49, 11, -37, 72, 3, 28, -66, -36, -48, 15, 15, 41, 3, 55, 55, -71, 49, -64, -37, -54, -6, 54, 1, -50, 8, -60, -44, -55, 28, -36, 61, -1, 50, -52, -5, -23, 51, 3, 14, -74, -60, -48, 42, 16, -69, 21, 18, 53, 30, 56, 75, -53, 32, -2, -28, -36, 13, 1, -16, -37, 38, -33, 38, 12, -10, -45, 62, -36, 31, -1, -35, 44, 26, -69, -16, 30, 25, 75, 6, -23, 53, 3, -1, 9, -75, 45, 46, 13, -30, -47, 52, -69, -5, 12, 16, 61, 42, 3, -51, -4, 75, -11, -36, 23, -7, 22, -25, -60, 21, 56, -8, -1, -17, 65, -70, -19, 34, 52, 70, -74, -71, 44, -68, -3, -20, 22, -18, -56, -53, 4, 13, -54, 66, 53, 42, -19, -3, -59, -4, -58, 73, 62, 14, -22, 49, 18, 35, 7, -6, 29, 6, -4, -5, 12, 68, 48, -42, -27, 65, -20, 52, 3, -1, 41, -22, -35, -54, 50, -19, 16, 65, -24, 0, 4, 30, -27, -56, -11, 53, 13, -60, -19, -69, 8, 68, 72, -20, -52, -31, -31, 1, -56, 45, 73, 60, -53, -38, -70, 72, 17, 19, 60, 66, -57, -14, 20, -9, 5, -69, -34, -60, -54, 23, -54, 27, 13, -58, -69, 37, -15, -26, -40, 4, -57, -42, -14, -36, -7, -11, -42, -68, -67, -58, 74, -49, 3, 16, 16, -68, 23, 57, -55, 42, 4, -36, -6, -58, -20, -2, 52, 40, 47, -64, -34, 64, -33, 27, -48, 36, -60, -15, 43, -52, 1, 39, -27, -74, -20, 62, -68, -73, 41, -48, 42, -32, -8, -40, -17, 47, 34, -41, 9, 3, -32, 50, -9, 9, 1, 18, -31, 14, -74, -66, 36, 0, 49, -67, 1, -47, 68, 8, -47, 33, 36, 70, -75, -50, -47, -19, 72, 60, 13, 5, -13, 57, -23, 54, -12, 53, -6, 32, -9, -7, 39, -49, 68, 12, -43, -8, 38, -51, 75, 64, 56, 33, 59, 54, 58, -66, -40, 52, 69, 48, -21, -20, 27, 31, -44, -61, 6, 26, 44, 71, -59, 8, -54, -66, -58, -23, -1, 54, -1, -2, 42, -21, -46, 23, -44, -66, 30, -9, 60, 23, -39, -37, -72, 62, 68, -41, 74, -2, 58, 43, -9, 75, -27, 13, -69, -12, 65, 5, -36, -12, -75, -71, 41, -46, 25, 72, -36, -20, -15, -52, -73, 19, -16, -72, 5, -26, -37, 4, 46, -57, -31, -39, -58, 15, 49, -52, -75, 36, 28, -35, -53, 29, -31, 61, 56, 69, 55, -56, -27, -36, -35, -26, 56, 23, -23, -14, 72, 13, 63, 42, 32, -46, -72, 47, 42, 50, 71, 42, 9, 21, -69, 29, -28, -27, 14, -47, -35, -7, -30, 11, 30, 9, 60, 10, -44, -40, 69, -50, 48, 56, 68, 2, -68, 69, -26, 49, 41, -31, 16, -26, 63, 20, -73, -40, 69, 14, -14, -42, -71, 29, 42, 34, -38, 27, -31, -9, 62, -38, 17, 32, -59, 7, -41, -54, 0, 8, 69, -37, 50, 9, 13, 37, -49, 13, 70, -58, -50, -22, -25, -46, -68, -60, 64, -31, 42, -45, 34, 26, -10, -25, -18, 4, 55, 16, 26, -21, -54, 17, 15, 71, -50, -50, 31, -26, 37, 25, -8, 62, -74, 40, -60, -67, 55, -74, -25, 21, -46, -67, -31, 20, -19, 27, -54, -40, -35, 45, 12, -13, -14, -48, -18, 9, -23, -65, 59, -62, 36, -25, 73, 37, -63, -64, 43, 68, -63, -58, 11, -35, -51, 56, 58, 5, 7, -72, 41, 47, 47, -23, -44, -43, 2, 12, 42, 55, 22, 23, 66, -20, 71, 64, -59, -68, 75, 57, 75, -66, 75, 9, -26, -54, -11, -44, 26, 69, -42, -11, 38, -71, 40, 70, -39, -34, 6, -75, -57, -48, 23, -66, 8, 16, 71, 22, 24, 70, 4, 21, -72, 1, -46, -22, 22, 18, 7, -30, 9, 40, 35, -28, 42, -3, -34, -72, 38, 45, -74, 55, 70, 23, 64, 2, -37, 57, -53, 60, 51, 24, 6, 54, -53, 33, -46, 44, -26, 35, -64, 58, -3, 44, -46, -36, -35, -7, -35, -74, -40, -34, 56, -45, 62, 42, 30, -50, 23, 52, -66, -2, 0, 13, -26, 22, -29, 2, -12, 20, -41, -2, 0, 31, -34, 28, 70, 7, -55, -43, 6, -21, -1, -14, 9, -17, -48, -37, 8, 48, -62, 16, -32, 13, -49, 15, -42, -5, -59, 19, -61, -27, -59, 13, -71, -17, -35, 72, 63, -17, -46, -7, 37, 26, 52, -30, -67, -74, 7, 15, 49, 20, -47, -59, -45, -21, 31, -14, 50, 46, -70, 62, -57, -56, -1, -55, 0, 39, -58, -13, -53, -31, 53, 57, 68, 29, -50, 74, 28, 32, 13, 1, -26, 39, 15, 2, -57, -31, 64, 66, -63, 69, 50, -45, -65, -26, -24, 11, -65, -9, 73, -45, 33, 49, -63, 25, 0, -38, 23, -47, 67, -41, 27, -35, 71, -33, 40, -62, 9, 28, -74, 21, 19, 52, 51, 30, -52, -51, -35, -44, 13, -40, -13, -32, -67, -3, 68, 9, 32, 14, 35, 21, 46, -14, 59, 41, 26, 23, 53, -41, -24, 52, 55, 70, 26, 29, 24, 49, 51, 62, -72, -13, -53, -12, 30, -45, 58, 23, 37, 14, -41, -6, -41, -73, 56, -58, 41, 4, 38, 18, 39, -62, -7, 16, -69, -57, -33, 28, 66, -57, 15, 69, 5, 37, -19, -43, 65, -37, 53, 25, 50, -64, -57, -69, -64, 72, -54, 53, 1, 59, -7, -38, 73, 61, 53, -74, -73, -57, 29, 68, -41, -32, 59, 37, -73, -38, 69, 68, 0, 47, 17, -28, 56, 33, -22, 68, 30, -3, 43, -45, -20, -40, -10, -25, -56, -33, -24, -54, -17, -70, -64, 17, -29, 70, -22, -26, -44, -28, -36, 29, -59, 54, 74, 72, 11, -26, 62, -35, 46, 29, -7, -52, 65, 58, -3, -69, -52, 48, -50, 6, 51, -39, -54, -53, -47, -1, -6, -18, 44, 33, -67, 60, 11, -69, 55, -56, -20, 41, -17, -52, -5, 51, -29, -18, 32, 41, -12, 55, 14, 11, -17, -13, 47, 4, 7, 73, -74, -75, -21, 45, 31, -13, 28, -34, -9, 7, -16, 44, -28, 42, 67, 42, 17, -40, -54, -29, -74, 7, -52, 13, -58, 7, 73, 62, -67, 5, 59, -66, 5, -40, 53, -41, 20, 3, -2, -67, -66, 57, 52, -21, 23, 41, -56, -37, 75, -35, 9, 74, 48, 33, 9, 63, -38, 6, 50, -30, -65, 31, -22, 14, 65, -47, 48, 7, 31, -30, 16, 40, -48, -10, -57, 48, -44, -38, -65, -47, 1, 18, -49, -29, -27, 35, -42, 10, -35, -68, 53, -26, 37, -45, 63, 24, -17, 35, -45, -62, -73, 46, 51, -48, -39, 68, -75, -10, -48, -67, 18, 28, 24, 42, 74, 72, 1, -43, 6, 39, -38, -16, -63, 72, 12, 73, 20, 71, 30, 51, -69, 33, 19, 56, 60, 55, 48, 58, -33, 75, 65, 60, 28, 13, 26, 24, 10, -51, 54, -62, 64, -61, -5, 74, -65, -68, 72, 31, -75, 26, 4, -69, -19, -53, 62, -36, -75, 32, -54, -33, 32, -67, -50, -18, 22, 49, -72, -46, 72, 58, -33, 58, 72, 38, 56, -69, 43, 50, 35, 43, -1, -37, 47, 55, -16, 32, -59, -16, -12, -37, 24, -56, -31, 47, -1, 66, 21, 3, -58, 15, -17, -15, -3, -21, -55, -23, -17, 63, -50, -59, 30, 24, -23, -1, 1, 36, -45, 18, -58, 19, 54, 40, 36, -53, 11, -42, -64, -46, 36, -47, 44, -59, 11, -35, -7, 31, 16, 51, 16, 41, 67, -32, -13, -33, 43, 63, -73, 73, 5, -55, 16, -19, 58, -25, 4, -7, 8, 15, 21, -34, 41, -11, -18, -23, 28, 50, -68, -34, 23, 24, -69, 13, 65, -9, 55, 32, -22, 55, 28, 57, 75, -34, -40, 55, 16, 39, -27, -52, -24, 67, -13, -58, -20, 44, -6, -70, 16, -1, -29, -36, -55, -25, 52, -65, 41, 29, 40, -58, 8, -8, 72, 6, 34, -44, -15, -26, 71, 31, -4, -31, 22, 58, -14, -75, 25, 53, -70, -35, -25, -25, 4, -5, 25, -22, 5, -11, -71, -30, 6, 13, 35, 2, -57, -7, 33, 1, 43, 26, -43, -39, 69, 54, -57, -21, 54, 43, -45, 58, -69, 5, -43, 8, 75, 55, 62, 3, -32, 66, 46, 49, 1, 5, -27, 19, 72, -71, -55, 37, 28, -25, 73, 21, -47, -62, 74, -70, 57, -47, 63, 63, 31, -58, -7, 30, 72, -21, -45, -35, -32, 74, -64, 44, 2, -15, -14, -2, -11, 4, -41, -59, 54, -46, 36, -71, -33, 34, -66, -54, 62, 70, -69, 17, -64, 0, -31, -67, 54, -2, -27, -56, -4, -16, 62, 71, 42, -30, -9, -47, 49, 23, -32, 25, 52, -72, 27, -56, 37, 35, -35, 21, 29, -28, -38, 39, 45, 4, 47, 21, -74, -58, 41, -4, -1, 25, -11, -36, 70, 56, -8, 41, 3, 35, -12, -22, 36, -61, -3, -3, 49, 35, -58, 1, -71, -23, -38, 49, 57, -69, -7, 56, -54, -42, -24, 20, 56, 39, 57, 50, 19, -26, 13, -56, -69, -75, -3, 41, -63, 67, -38, 60, 25, -22, -15, 29, 30, 22, 1, 9, 26, 69, -10, 47, -51, 39, -11, -71, 2, -29, 52, -57, 18, -11, -37, 24, -11, 35, -11, -1, 25, 25, -17, -26, -75, 43, -75, 30, -13, 1, -38, -63, -8, 27, 57, 14, -12, -29, 16, 66, 17, -8, -67, -41, 54, -31, 56, -35, -71, -32, 40, 29, 66, -53, -75, 66, 64, -75, 18, -25, 0, 55, -14, 67, 6, -33, 4, 70, 11, -56, 58, -48, 10, 64, -16, -12, -42, -35, 29, -38, 6, -7, 64, -4, 13, 64, -16, 1, 64, -74, 50, -12, 57, -42, -22, -15, 0, 55, -23, -66, 74, -41, -39, 6, -52, 21, 70, -19, 59, 21, 16, -13, -64, 2, 56, 24, -10, -36, -50, -24, -35, 73, 38, -56, -45, -62, 5, 28, 68, 57, 37, 64, -61, 74, -5, -38, 17, -13, 16, -2, -68, -46, 60, -57, 31, 40, 40, -57, -74, 63, -8, -36, 60, -46, -16, -61, -35, 62, 41, -45, 43, 2, -58, 55, -2, 12, -61, -61, 74, 30, 10, -72, 59, -8, -56, 14, -44, 59, 30, -45, 47, -53, -5, 29, -26, 54, 42, 15, 40, 7, 43, 5, -67, 60, -17, 7, -6, -3, 19, -10, -50, -48, -7, -67, 19, 12, 21, 49, -6, -25, -72, -37, -3, -2, 67, 47, -26, 31, -16, -64, -38, -49, 15, -31, -66, 73, 51, 3, -6, -8, 69, 19, 19, -16, 26, -37, 70, -31, -66, -12, 17, -63, 24, -63, 9, 13, 59, 58, -31, -35, 68, 6, -11, 7, 48, -2, 4, 21, 75, 71, -62, 68, 13, 30, -24, -39, 66, -32, 5, 75, 31, -54, -65, -21, -42, 19, 68, -61, -1, -41, -23, -9, 38, 42, 73, 11, -38, -1, -44, -39, -7, -33, -49, -70, 73, 1, -36, 61, 44, 44, 59, 0, 63, 69, 52, -54, 12, 42, -42, -67, 74, 11, 0, 37, -25, -5, -28, 12, 68, 1, 47, -15, 44, 73, -12, 39, -2, 27, 22, -33, -7, 5, 40, -20, -2, 14, -1, -68, -21, 33, -59, -23, -34, 14, -62, 16, -67, -17, -50, 74, 60, 72, -19, 26, 70, 44, -13, -10, -7, -67, 32, 59, 14, -6, -36, -66, -69, 36, -58, -15, -7, -44, 37, 32, 45, 49, -28, 51, -44, -2, 50, -62, -6, -45, 39, -14, 73, -52, 52, -12, -43, 6, -28, 46, 74, 9, 55, -71, -31, 70, -11, 36, -50, -52, -8, 70, 72, 38, 46, -49, -42, 20, -36, 25, 48, -74, -66, 45, -51, 61, -42, -19, -11, 3, -51, -15, -64, -73, -11, -22, 72, 51, -64, -53, 75, 2, -61, 71, -38, 60, -54, -5, 2, -16, -56, -25, -15, -47, -58, 7, -64, -25, 62, -1, 53, -65, 59, 62, -63, -29, -37, -68, -54, -26, -46, -55, 49, -32, -61, -65, -49, -42, 5, 26, 15, 23, -75, 73, 49, -57, 5, 59, -9, -11, -18, -33, -1, -35, -47, 10, 11, -9, 17, 31, 39, 44, 49, 12, -66, 63, 23, -40, -56, -48, 62, 32, 48, 60, 30, 22, -73, -43, 5, -8, 21, 60, 34, -58, -51, 62, 27, 34, -24, -34, -13, -61, -66, -40, 26, -56, -54, -29, -23, -35, -1, -37, 70, -31, -52, 24, 66, -52, 56, -7, 13, 1, -23, -29, 19, 0, -42, -32, -44, 7, 10, 18, 21, 17, 53, -31, 34, 74, 16, -64, -39, -63, -28, -44, -19, -7, 53, -30, 15, 32, 38, -48, -45, -62, -1, 47, 11, 30, -60, 42, -39, 23, -18, 55, -38, -41, -54, 72, -44, 37, -68, -10, 47, -23, 19, -47, 46, -3, -4, -15, -47, -44, 12, -19, -31, -65, -47, 55, 38, -32, 19, 74, 64, -75, 51, -50, -42, 73, -54, -11, 34, -49, 52, 4, 2, -4, 32, -28, 66, -50, 32, -59, -19, -34, -3, 24, -25, 25, 3, -63, 66, -55, -66, 54, -55, 60, -73, -24, 57, -54, 38, 14, -29, 15, -58, 48, -65, 47, -56, 74, 72, 49, -61, -25, -63, 11, 74, -13, -41, 0, 0, -51, 20, 9, -74, 38, -7, -72, -61, -27, -51, 52, 60, -5, -9, -74, -35, -1, 46, -16, -5, 40, -45, 9, -61, -32, -57, -62, 30, -25, 13, -48, -1, -45, 34, -2, 68, -48, 1, -69, -2, 24, 57, -18, -59, -30, -19, -18, 45, -49, 41, -38, 66, 70, 47, -73, -38, 63, -60, 65, -38, 26, -58, 34, 56, 51, -43, 47, -75, 31, 51, -4, -21, 32, 53, -4, -73, -44, 53, 45, -18, 16, -69, -30, 8, 51, -29, 43, 36, -16, 33, 73, -65, 48, 30, 64, 21, 62, 35, 20, 15, 9, -60, 70, -35, 67, -12, -35, -53, -37, -68, 3, 52, -63, 46, -15, 61, -59, -48, 22, -1, 58, 17, 9, 28, -29, -5, -26, -45, -47, 67, 46, 37, -71, 38, -74, 71, -52, -35, -59, -14, -30, 17, -40, -18, -15, 20, -32, 0, 46, 65, 74, 28, 4, 5, -19, 51, 75, 28, -70, -48, 19, 49, 64, 23, 11, 64, 17, 34, -49, 31, -58, -4, -28, -22, 54, 32, 71, -56, -44, 41, -69, -48, -8, 10, 32, 46, -15, 32, -4, -11, 57, -63, -38, 44, 35, 47, 30, -26, 3, 56, -71, 21, -24, -24, 72, -48, -69, 67, -29, -40, 31, -25, -12, -53, 61, -56, 66, -32, 49, -14, 30, 29, -2, 66, -3, -45, 35, -49, 3, -38, -69, 7, 56, -20, 57, 52, 8, 61, 42, 52, -55, -3, -50, 6, 17, -67, 24, 7, -24, -3, 66, -71, -52, -14, 70, 20, 14, 29, 44, -59, 64, 48, 22, 43, -47, 3, 19, 34, -14, -17, 8, 6, 55, 33, -65, -6, 41, 34, -75, -60, -47, 64, -58, -23, -28, -64, 70, 62, 38, 39, -75, 24, 9, 22, -9, 37, -53, -67, -7, 8, -9, 75, -63, -31, 32, -53, 38, -4, 56, 37, 9, -69, 25, 26, -17, 71, 35, -24, 55, -5, -61, 55, -59, 21, 2, 8, -19, 22, 14, 49, -45, -71, 48, -33, -27, 3, -11, -66, 72, -33, 46, 3, -27, -7, -49, 30, -12, 59, -70, -33, -24, -58, -53, -8, 38, 22, 73, -57, -32, 11, 66, -4, 14, 38, 38, 60, -37, -51, 69, -43, -9, 39, 35, 38, -43, 61, -8, 20, 42, -3, 61, -58, 12, -68, 10, -26, 27, 7, -7, 68, -59, -17, -11, 30, -57, -51, 14, -20, -26, 8, 12, 38, -29, -30, 0, 1, -47, 65, -54, 71, -14, -69, -63, 73, -64, 22, -30, 36, -48, 36, 28, -32, -59, -59, 73, -41, -34, 9, 12, 13, -59, -51, -25, -14, -6, 51, 62, 20, 40, -70, 15, -51, -66, 28, -56, -55, -26, -11, 56, 1, -51, 7, 42, -35, 23, 39, -2, 62, -27, -66, -1, -13, -44, 50, 48, 23, 23, 33, -32, -15, 38, 58, 7, 48, 10, 27, 66, 58, -62, 45, -19, -39, -24, -52, -1, 72, 60, 70, 59, -45, -71, -20, 18, -42, -48, -12, 55, 50, -55, -55, -42, 59, -73, 38, 29, 11, -13, 19, -9, 1, -12, 47, 35, 39, 68, -42, 36, 51, -47, 17, -70, -45, 72, 21, -14, -51, -66, -35, 72, -48, -15, -48, -65, -14, 66, 37, 70, -23, -19, -15, 51, 44, -46, 10, 6, -55, 42, -36, 71, 68, 56, -75, -55, 50, 22, 6, 74, 29, 45, 69, 56, -46, -55, 65, 13, -65, 26, 7, -14, -69, 65, -41, 49, -58, 43, -23, -38, 9, 16, -43, -1, -6, -45, 19, -32, 50, -51, -35, 1, 69, -42, -18, -54, -24, -31, 34, -13, 70, -36, 46, 75, -49, -71, 46, -32, 47, -53, 3, -22, 36, 33, 52, -48, 64, -5, -7, 36, 20, 33, -38, 11, 64, 17, 32, -35, 59, -11, 25, 53, 28, -7, 50, 54, -3, 20, -55, -33, 40, 23, 18, -2, -19, -5, 25, -31, 65, -59, -73, 7, 49, -38, -57, 36, 52, 48, 74, 35, -39, 21, 11, 62, -62, -15, 41, 8, -72, 61, 48, 41, 6, -9, -36, 62, 61, 62, -47, 48, -73, -44, -22, 50, -9, -6, 8, -32, -34, 6, -75, 1, -49, 9, -13, -36, 68, -50, 45, 71, -67, 18, 34, 15, -67, 71, 1, 67, 58, 28, 37, 58, 57, -61, 32, -28, 6, -36, 13, 46, 45, 12, -29, 69, -55, 31, -45, -63, 57, -75, -70, 65, 16, 40, 2, 22, 35, -74, 13, 15, 29, -26, -2, 10, -13, -46, 55, 68, -8, -7, 36, -41, -73, -69, -47, -53, 38, -19, -42, 19, -21, -37, 6, 70, -75, -69, 16, 36, -68, -49, -27, 36, -1, 46, -32, 61, 74, -53, 51, -10, 13, 12, 24, 15, 16, 50, 38, -22, -44, 71, 70, 10, -44, -1, 3, -43, 5, -57, 66, 12, -30, -37, -30, 44, -66, 13, 27, -70, 35, 0, -5, -27, -66, -59, 63, 26, 65, 23, -74, -57, 16, 72, 26, 48, -7, -47, -71, 73, -30, 70, 7, 13, -45, 52, -21, -38, -13, -70, -33, -54, 3, 35, -8, 13, 50, -22, -37, 39, -75, -36, 57, 17, -42, 7, -11, 24, 34, -9, 19, -72, -17, -50, 16, 13, 75, 70, 49, -16, 73, -60, 6, -2, 49, 71, -65, 23, -27, -29, -14, -26, 9, -35, 64, 42, 45, -25, -11, 3, 41, -68, 4, -52, -44, -56, 34, -47, -64, 5, 13, -69, 21, -59, 5, -8, -64, 13, -61, -15, 60, -2, 32, -7, 36, 20, -43, 5, 68, 21, -69, 33, 29, 10, 54, 60, 28, 10, -63, 37, -60, 25, 42, 34, 39, -29, -50, 51, 57, -38, -42, 41, 35, 65, -42, -5, 7, -9, 73, -1, -64, -72, -46, 38, 12, -70, 22, -38, 15, 33, 74, 28, -20, 38, -14, -56, -67, 9, 70, 66, 46, -50, 29, 3, -63, 63, 71, 17, -24, 69, -60, -15, 70, -33, -52, 4, -30, 43, 41, 60, 0, 38, 13, 54, 0, 72, 73, 7, 6, 65, -5, -24, -61, -52, 55, -51, -67, 50, 41, -16, 41, 54, 43, 34, -55, 66, -38, -10, 31, -72, -28, -44, 39, 58, -66, -37, 53, -71, 43, -17, 67, -38, 32, -70, -16, 9, -46, -8, -18, 70, 50, -55, 46, 17, 54, 66, 5, -59, -22, -40, -58, 23, -11, 56, 6, -4, -59, -17, 0, 58, 39, -9, -56, -5, -6, 1, -73, 21, 69, -16, 13, 41, 4, -17, -18, -19, -29, 60, -3, 24, -56, 12, -28, 9, -10, 51, -71, 6, -44, 3, -14, 70, 69, 6, -13, -14, -69, -11, -69, 73, 46, 18, 38, -27, -75, -58, 29, -28, -74, -52, 69, -56, 35, -37, 26, -51, -62, 28, 28, -31, -45, -61, -37, -53, 18, 24, 6, 22, -63, 12, 18, 59, -46, -20, -46, -47, -4, 58, 0, -5, -72, -9, 14, 38, 30, -38, 60, 43, 66, 12, -65, -57, 24, -29, -37, -36, 70, 44, 60, -68, -21, 2, 64, 6, 55, -60, 32, -25, 73, -46, 46, -75, 21, -18, 36, -25, 20, 20, -60, 8, -46, -52, 24, 52, -5, 63, -62, -11, 29, 73, -6, -70, -1, -20, 12, -21, -5, -32, 27, -10, -2, -5, -12, -59, 53, -54, -11, -5, 39, 4, -73, 69, 28, 26, 43, -55, 11, 56, 7, -35, 54, 75, -32, -25, -21, 55, 27, 48, -54, -21, -40, 17, 49, 22, 31, 24, 43, -56, -57, 7, 21, -57, -2, -29, 43, -35, -9, -22, -55, 74, 16, 72, 71, 60, -28, -28, 37, 74, -56, 56, -25, -22, -5, -51, 75, -50, 48, 42, -31, 65, -29, 66, -68, 44, -39, 50, -67, 26, -49, -48, 22, 42, -54, 17, 24, -9, 64, -14, -10, -69, -36, 38, -18, 35, 62, -19, 58, 33, -55, -48, 20, -8, -60, 27, -42, -26, 0, -35, 75, 26, -10, 19, -10, 11, -40, -61, -73, -53, -2, -10, -49, 35, -48, 8, -6, -63, 62, -25, 43, -69, 0, -13, -4, 15, -64, 28, 62, 11, 68, 60, -41, -18, 3, 25, 68, 37, 37, 68, 59, -43, -18, -66, 67, 10, 15, -16, 20, 1, 34, -13, 5, -42, 47, -74, 46, 58, 29, 32, -6, 19, 16, 26, -75, -58, -25, 68, 54, -66, 61, 37, -34, -35, 44, -44, 48, -17, 15, -8, 57, -27, 52, -14, 4, 23, -13, -26, 6, -62, -72, 73, 32, 18, 23, 30, 35, 72, 21, 13, -70, 4, -28, -30, 44, -62, 1, 17, -4, -60, -69, -23, -14, 59, 36, 65, 6, -54, -39, -66, -41, -36, -69, 65, 55, 30, 19, 14, 24, -38, -51, 29, 41, -6, 74, 10, 7, -1, -49, -75, 12, -45, -25, 73, -62, -64, 60, 18, -43, -57, 27, -11, -19, 34, -22, -40, -14, 71, 48, -66, -43, 72, 36, 74, -9, 33, 6, 71, -44, 30, 72, 42, 60, -29, 39, 74, -18, 22, 16, 12, 40, -35, -74, -55, 74, -23, -21, -18, -30, -49, -11, 1, -55, -50, -3, 9, 58, -73, 5, -64, 32, -1, 53, 14, 45, 15, 12, -50, -41, -50, 35, 74, -9, 36, -58, -13, -64, -6, 43, -19, 20, -44, 55, 38, -21, -24, -28, -41, -24, 50, -29, -68, -27, -54, 20, -60, 36, -44, -37, 68, -20, 74, 67, 44, 32, -69, -47, 43, 0, 71, -53, -58, -50, -74, 55, 2, -24, -51, 37, 27, 72, -70, 33, -31, -49, -23, -17, 61, 6, 21, 53, 59, 17, 42, 27, -26, 48, 54, -61, -30, 47, -41, -13, 72, -41, -35, -3, 8, -13, -42, -41, -16, -37, 67, 26, -11, -34, -67, -28, 48, 28, -50, 31, -31, 65, -19, 16, 38, -43, 29, -70, -72, 61, -9, 74, -56, 31, -5, 27, -60, 28, 60, -1, 64, 49, -50, -25, -60, -44, 23, 61, 59, 46, 14, -49, 35, 68, 40, -5, -51, -7, 1, -47, -21, 67, -51, -4, 20, 19, -54, 33, -31, -70, -43, -43, 54, -20, 7, 67, 11, -48, 52, -7, 73, -9, 19, 31, -17, -17, -50, 8, 50, 24, 34, -49, 13, 56, 20, -43, -1, 41, 66, 41, 46, -55, 71, 23, 0, 2, 14, -67, 28, -11, 1, 23, 55, -58, -22, -40, -1, 4, 41, -29, -50, -1, -3, 39, -21, -59, 71, 51, 58, 59, 16, 26, -74, 11, -29, -1, -64, 61, 8, 37, -26, -69, -16, -49, -53, 38, -14, 21, -36, -48, 67, -11, 24, -14, -48, -74, 0, -54, 50, -20, -73, -9, -69, -73, 75, -25, 1, -67, -42, -69, 43, 5, -64, -48, 31, -42, 63, -60, 52, -51, -35, 41, 11, 64, -51, 37, 63, 24, 56, 38, -71, 56, -49, -67, 58, -52, -17, -18, -45, 17, -14, 73, -56, -3, -53, 51, 28, -68, 64, 2, -44, -47, -35, 41, -61, -11, 2, -75, -62, -20, 38, -60, -40, 64, -52, -59, -66, 4, -2, -36, -57, 57, -38, -37, -23, -16, -64, -71, -10, 75, 5, 21, -50, 43, -14, -38, -43, 61, -38, -32, -35, 75, -17, 1, 61, 6, 17, 71, -68, -63, -41, -49, 69, -6, -11, -30, 52, 0, -27, -34, -3, 51, 62, 22, 18, -29, 59, 50, -46, -54, -58, -5, -57, -2, 69, -71, -74, 8, 75, -66, 20, -42, -40, 11, 28, 24, 57, 4, -54, -48, 45, 18, -73, 29, -36, 20, 73, -55, -7, -48, -36, 8, 22, -17, -69, 15, -13, -68, -55, -14, -59, 40, 17, -24, -25, -33, 73, -46, 44, -57, -21, 11, 36, -19, -35, 73, 75, -38, -59, -8, -13, -20, 73, -67, 38, -72, 21, -51, -66, 41, 8, -50, 3, -50, 0, 52, -10, -3, -72, -41, 14, -17, 45, -26, 37, -68, -30, 36, -32, -14, -50, 30, 41, -52, 37, 2, -49, -18, 26, -40, -54, -43, -16, 22, -20, 59, -2, 45, -22, 0, -72, 67, 58, 47, -36, 19, 54, 7, -22, -54, 68, 3, 50, 31, 24, 11, -43, 51, 66, 57, -67, -64, -62, -10, 32, -7, -29, -48, -38, 25, 27, -36, 14, 7, -67, 51, -51, 60, -18, 2, -69, -28, -73, 54, -72, 27, -11, -42, 0, -21, -61, 6, -11, -50, 72, -55, 18, -35, -28, 54, 63, 73, -60, 2, 4, -52, -25, 28, -68, 33, -48, -64, -73, -47, 65, -70, 55, -22, -38, -23, 31, -24, 58, -56, 0, 52, -36, -58, -58, 9, 69, -71, 6, -67, 4, -65, -46, 55, 36, -38, 10, 62, -29, 12, -61, -39, 16, 67, 12, 53, -34, -33, -49, -52, -14, 26, 74, 23, 42, -60, -43, 35, -58, 38, 44, 22, 46, 73, -1, 7, -43, -67, -9, 4, 20, 3, 38, -40, -8, -26, -65, 33, 15, -38, 54, -75, 63, 52, 22, 27, 65, 54, -13, -70, 16, -45, 27, -15, -50, -52, 65, -17, -44, -20, 60, 49, 58, 22, -66, -28, 69, -58, -71, 8, -21, 56, 7, -35, 31, -47, 67, 18, -71, -22, 23, 18, 6, -28, -73, 30, -5, 67, -65, 26, -29, 70, -2, -49, 14, 5, -2, 5, 22, 0, -62, -74, -19, 18, -36, -66, 44, -47, 27, 48, 7, -25, -10, -65, 22, -9, 38, -60, -18, 48, 41, 27, 40, -39, 51, -22, 41, -26, 57, -12, 47, 70, -13, -50, 10, 26, -41, -22, 54, 62, -50, -17, -41, 13, -8, 56, -72, -46, 71, -16, -73, 35, -65, 40, 71, 61, -59, 35, -43, 73, -53, -71, 67, 7, -48, -1, -43, -13, 52, -67, -29, 75, -10, 5, 12, 55, -15, 14, -67, -21, 73, -67, -64, -68, 49, -71, 66, 65, 39, -52, 60, 61, -50, 49, -10, -23, -28, 22, 37, -52, 29, -68, -53, -59, 12, 32, 71, 71, -30, -72, -26, -33, -65, -15, -28, 57, -13, -39, 44, -49, -18, 28, -66, 7, 1, 0, 57, 48, -56, 19, 69, 46, 26, -60, 62, -37, 45, 57, -42, -60, 59, 5, -20, 67, 63, 26, 48, -26, 62, 16, 0, -32, -34, 8, 48, 42, -68, 29, 12, -49, -28, 5, 71, 72, 18, 57, -41, -13, 37, -10, 0, 20, 70, 56, 11, 55, 6, -19, -47, -10, 70, 27, 33, -40, -41, 5, 75, -36, -44, 9, -12, 2, -62, -17, -2, 29, -35, 30, -62, -74, -58, 14, 19, -66, -6, -48, 64, 73, 6, -61, -13, 0, 41, -58, 33, 73, 22, 32, -39, 51, -35, 23, -23, -24, -70, 48, -73, -32, 2, -60, -33, 19, 29, 59, 28, -55, -65, 14, -60, 14, 29, 2, -62, -6, 19, 46, -10, -37, 0, 24, -63, 38, -29, -11, -64, -25, -38, -62, 18, 37, -48, 59, -19, 56, 42, -69, 75, 51, 19, -61, -11, -28, 15, 1, 39, -44, -31, -47, -7, 45, 53, 5, 5, -54, 69, 17, -4, -47, 30, -63, 66, 55, 71, -31, 36, 35, -27, 33, 10, 67, 45, 73, -37, -16, -4, -73, 16, 40, -47, -67, 7, -70, 11, -63, -48, 4, 29, 21, 31, -19, 33, 21, -39, 28, 65, 70, -14, -38, 25, 71, -46, -6, 66, -10, 54, -14, -10, -8, -51, 19, -2, 31, 22, -67, 43, 47, 10, -6, -7, -35, 51, -50, 61, -66, 52, 48, -74, -38, -67, 26, -45, -40, -56, -56, 25, 71, 5, -60, -13, 27, 34, 58, -17, -20, 66, -50, -50, -1, 20, 18, 39, -7, 41, 23, 0, 17, -7, 1, 52, 1, -51, -68, 36, -32, -51, -16, -36, 29, -1, 26, -21, -45, 9, 37, 8, -3, 62, 33, 71, 4, -25, 33, 70, -59, -22, -8, 31, 46, 66, 8, -28, -61, 13, -70, -17, 37, -11, 20, -12, 61, -30, 42, -60, 52, 3, 22, -28, -12, -21, -35, 65, 28, 73, 58, 42, -27, -26, -3, -56, -35, -73, -9, -23, 13, -4, 35, -26, 59, -21, 38, 44, 23, 2, 60, -3, -70, 6, 42, -9, 58, -68, -22, 8, -73, -40, -26, -24, 8, 45, -5, 46, 45, 59, -53, -17, -23, 58, 32, -40, -41, -8, -71, 55, 70, 62, -23, 73, -10, -59, -14, -30, -54, 39, 54, -51, 75, -48, -2, 5, 70, 66, -25, 40, 47, -3, -53, -52, -23, 54, -18, 10, -31, -16, -11, -39, -32, 39, -42, 33, 56, 19, -73, -74, -20, 56, -52, -23, -69, 19, 57, -75, 9, -44, 40, -20, 27, 60, 2, -72, 37, 57, 13, -70, -35, -73, -34, 6, 39, -3, -37, 17, -62, -37, 19, -7, -58, 40, 44, -54, -16, 25, -56, 66, 55, 58, -31, 6, 42, 46, 7, 3, 25, -55, 6, 65, -55, 45, -7, 59, -34, 29, -1, -23, 67, -58, 44, -69, 57, 12, -50, -37, -41, -30, -46, -62, -48, -2, 19, 69, -34, -49, -5, 66, -31, 74, 53, -13, 44, -30, -32, -68, 74, 42, -17, 63, 59, -49, 68, 39, 36, -58, 75, 70, -13, -47, -67, 12, 24, 25, 4, 65, 49, 72, 53, -60, 70, 30, 2, 36, 73, 46, 44, 69, 12, -49, 57, -6, -25, 49, -45, -65, 64, -46, -71, -26, -19, -65, 61, -73, 36, -11, 66, 7, -15, 43, 23, -20, -4, -51, -62, -9, 70, 57, -15, 5, -70, -34, 72, -20, -63, -49, -10, -75, -22, -7, -26, 32, 3, -42, 35, -37, 22, 25, 44, -70, -10, -9, -17, 59, 15, -4, -25, 8, -24, 35, -65, -19, 74, -69, 35, -65, -43, -53, -67, 8, 15, -19, -35, -57, 14, 75, -21, -42, 22, -53, -37, -64, 13, 21, 69, -49, -60, -32, 34, -9, -73, 44, 47, -75, 48, 6, -67, -71, 29, -61, 10, -34, -5, 50, -16, -69, 47, 37, -35, -7, 59, 3, 3, -5, -53, -4, 21, -38, 37, -23, 26, 39, -57, -3, 37, 66, -74, 43, 68, 28, 57, 2, 69, -25, -25, -24, -19, -54, -63, 21, 13, 71, -53, -62, -12, -33, 7, -67, 2, -32, -17, -48, -71, -1, 22, 39, -11, 21, 4, -21, -27, -15, 55, -33, 33, -46, 18, -61, -27, 30, 33, 59, 23, 53, 70, -64, -58, -1, -58, 19, 40, -1, 44, 42, 73, -11, 5, -13, -66, -69, 39, -17, -10, 18, 23, -53, 45, -37, -39, -59, 66, 68, 75, 11, 45, 68, 20, 63, -9, 38, 4, -44, -39, -29, 73, -42, 35, 1, 18, 44, 7, -20, -51, 72, 73, 47, -56, 41, -68, -22, 57, 71, -32, 54, 7, -62, 46, -49, 74, -40, 62, 0, -9, -53, 46, -12, -21, 5, 62, 70, -28, -6, -26, -4, -10, -30, -34, 7, -67, -29, 61, 63, -33, -47, 41, 49, -36, 10, 75, -40, 45, 60, 34, -40, -69, 4, 21, -17, -68, 8, -24, -21, 75, 23, 48, -11, 68, -64, 72, 74, -17, 55, 61, 25, -70, 25, -2, -32, -41, -5, 1, -74, -21, -41, -41, -16, 39, 55, 40, 44, -15, -62, -53, -16, 37, 68, 47, 27, -71, 41, 26, -13, 18, 11, -66, 23, -40, 5, 64, -8, 73, -10, -7, -25, 24, 27, 34, -13, 5, -4, -47, 65, 10, -27, -28, -29, -34, -57, 73, -32, 57, 21, 30, -1, -45, 37, -54, -10, -34, -65, 56, -37, -2, -27, 13, -54, 74, -31, 7, 3, 41, 35, -10, -27, -67, 37, 17, -26, 53, 12, 17, 34, -42, -31, -43, -12, -70, -23, 51, -31, -15, 29, 7, 58, -75, -55, -72, 74, -11, 10, -1, -48, -32, 64, -2, -24, 24, -61, 23, -1, 25, -38, -44, 56, 6, -12, -32, 9, 38, -59, 53, -53, 46, -18, -73, 46, 2, -69, 42, 65, 14, -35, -61, 57, -49, 11, -45, 50, 23, 53, -28, -28, -61, 3, -48, 18, 64, -7, -49, 25, 8, -74, 47, -22, -16, 48, -54, 59, 52, 63, 46, -10, -48, 59, -30, -22, -8, 0, -49, -61, -22, -4, -15, -10, 74, 12, -67, 60, -72, -43, 9, 11, -41, -21, 64, 16, -49, -68, -3, -73, 70, -34, -10, -54, -53, 35, -3, 14, -42, 21, 28, 9, -59, -63, 74, -61, 23, -69, 75, 26, -36, 6, -39, -4, 60, -53, -66, -67, -46, 6, -65, -52, 45, -1, -33, 67, -44, 37, 5, -11, -17, -44, 73, -1, -32, 72, 14, 66, -75, 11, 14, -36, -61, 48, 33, 75, 70, 42, -70, -54, -29, -59, -33, -60, 13, 7, -70, 44, -31, 8, -42, 27, 39, -47, -50, -68, -51, 37, 71, -52, -30, 8, -13, -17, -20, -55, -20, -25, 60, -15, -6, -45, -1, 37, -31, -64, -32, -26, 56, 10, 55, -64, -39, 19, -36, -15, 24, -13, -56, 19, 10, -10, -49, 70, 46, 7, -63, -50, 55, 73, 10, -29, -50, -66, -70, -8, -55, -28, 39, 74, 57, 19, -66, -59, -38, -28, 1, 61, 32, 20, 2, -34, -68, 27, -42, 53, -42, -29, -73, -65, -34, 11, -21, -9, 20, -15, 59, 38, 32, 22, 35, 13, -35, 44, 27, 0, -62, -48, -15, 45, 46, 61, -67, 51, 12, -33, 27, 45, 11, 29, 53, 52, -38, -46, -35, 57, 14, -52, 18, -30, 44, -23, 57, -69, -57, 8, 7, -43, 34, 65, 75, 2, 50, -67, -23, -14, -27, -72, -47, 59, 31, -72, 33, 68, -42, 73, 48, 47, -56, -10, -60, 63, 42, 70, 67, 60, 0, -4, -61, -44, -16, -61, 33, -42, -55, -67, 18, -7, -64, 44, -26, 40, 48, -69, 31, -72, -72, 3, 48, -53, 68, 61, -68, 32, 53, 75, 16, -22, -7, 31, 7, 52, 43, -35, -67, 63, -29, 26, -22, -18, -8, 27, -55, -38, 31, 51, -35, 34, -22, -64, 57, -32, 72, 62, 75, 50, 61, 15, -50, -21, -32, 32, -45, -67, 70, -39, 69, -35, 62, -29, 21, -23, 71, 39, 14, 26, 14, 55, -15, 67, 66, -36, -43, 60, -50, -44, 32, -66, 44, 57, -14, -63, 12, 14, -57, 4, 51, -63, 43, 35, -17, -14, -64, -21, -51, 26, -73, 38, 3, -13, 27, -9, 24, 59, -25, 50, -61, -68, 57, 58, 62, -33, 68, -2, 56, -64, -73, 29, -52, 43, -11, 4, -47, 0, 56, -23, -50, 59, -61, 26, -30, 39, -59, 68, 22, -10, 42, 36, -3, 21, 16, -17, 63, 9, 55, 41, 18, 55, -5, 39, 22, 57, -33, 50, -19, -52, -51, 5, -69, -39, -45, -26, 75, -28, -34, 21, 35, -70, -21, -44, 24, 70, 12, 11, 1, -11, -25, -59, -32, 43, 55, 63, 24, -55, 35, -73, -32, 59, 7, -28, -56, 36, 19, -59, -70, 59, 37, 40, 64, -60, 71, 13, -67, 5, -54, 7, 70, -6, 24, -40, -41, 1, -52, 58, 21, 56, 61, 62, 38, -10, -44, 55, -50, 51, 72, -45, 32, 33, 70, 18, 47, 63, -47, 53, -7, -27, -16, -15, 42, -70, 20, -74, 7, 41, 57, -50, 22, 42, -63, -18, -43, -34, -39, -20, -61, -43, 11, 46, 64, 5, -11, 33, -7, 17, 10, 59, 65, 67, -32, 30, 73, 63, 31, 4, 27, 10, 27, -29, -25, 37, 28, 5, -72, 64, 60, -58, -56, -5, 62, -70, 74, -25, 36, -11, 65, -30, -28, 55, -39, 13, 7, -44, 0, -40, 33, -51, 45, -15, -5, -56, -54, -53, 24, -51, -66, 9, -35, -49, -74, -49, -44, 75, -1, 67, -12, -12, -41, 33, -35, -7, -30, 47, 25, 44, -69, -18, 68, 50, 42, -12, 69, 62, 8, 16, -65, 17, -53, -27, 43, -52, -1, 72, -52, 71, 61, 9, -16, -56, -35, 22, 13, 10, -8, -38, -24, -4, 17, -31, -30, -18, 30, -38, -32, -38, 53, -24, 53, 75, 25, 18, -55, -54, 15, -32, -58, 0, 51, -1, 20, -60, -55, -45, 25, 12, -10, 75, -69, -69, -32, -24, -12, 71, 13, 31, -43, -12, -68, -68, -15, 30, 26, 6, 51, -35, 47, 66, 38, 22, -11, -20, 35, 8, 10, -17, -58, 73, -18, -52, -71, 25, 0, -10, 20, -65, -56, 50, -3, -51, 58, 57, 54, 8, -15, 27, 46, -43, 18, 8, 52, -71, 64, 12, 12, -4, 70, 30, -6, -24, 53, -2, 74, -25, 61, 16, -16, -73, -12, 56, -49, -30, 35, -73, 51, -57, 28, 19, -25, -30, -48, -51, -28, -62, 36, 60, 9, 28, 12, -73, -74, -13, -2, 75, 36, -18, 13, -56, -16, -74, 73, 9, -31, 30, 11, -57, 48, -37, 37, -55, 6, 62, -30, 54, 73, -72, 36, 7, 32, -30, 7, 33, 32, -72, 31, -8, -15, -32, 9, 42, -33, 6, -25, 12, -39, 60, 28, -67, -53, -11, -46, 27, -26, -3, 3, -29, 0, -37, 51, -46, 8, -19, 63, -38, -18, 16, 28, 40, 57, -39, 6, -51, 41, 55, 34, -74, 39, -14, -68, 61, 48, -41, 10, -54, 31, -63, -9, -44, -25, -36, -15, 56, 20, -30, -57, -74, 59, 44, 39, 41, -71, -30, 63, 45, -51, 21, 44, 63, -69, 52, 46, 54, -65, -21, 74, 40, -9, -11, 69, 40, 26, -24, 18, -29, 20, 34, -30, 3, 2, -66, -34, 7, -23, -47, -24, -1, 47, -57, -16, 53, 70, -48, 30, -73, 6, 26, 40, 71, -63, 33, 35, 38, -68, -23, -69, 27, -64, -25, -48, 13, -18, -6, -58, 34, 22, -8, -45, -8, 10, 14, -31, 2, 41, 72, 4, -30, 20, -31, -35, 32, 75, 75, -5, -69, -26, 1, 33, -17, 49, 61, 70, -45, -23, -64, 62, 72, 3, -59, -12, -65, 30, 31, 12, -6, 27, -59, 39, -28, -17, -74, -74, -20, -75, -4, -13, -28, 71, -58, 31, 44, -75, 25, 75, -23, 34, 61, -26, -40, -73, 37, -30, 30, -8, 58, -54, -58, 72, 58, -13, -23, 59, -12, 32, 57, 60, -57, -46, 53, -41, 58, 19, -41, 7, 18, 12, -37, 2, 61, -2, 2, 20, 44, -46, -63, 26, -24, -48, 20, -44, 14, 72, -60, -74, 28, 72, 59, 45, -52, 34, -72, -70, -22, -38, 10, 69, 47, 49, -5, 32, -29, 70, -25, -61, -51, -13, 38, -2, 14, -18, 29, -50, -24, 44, -49, -71, 39, -67, 47, 62, 42, 48, 68, -56, -66, 2, -62, 57, -25, 6, 11, 20, 1, 61, 34, 23, -30, -5, -57, 57, 52, 47, -69, -49, 14, -44, -47, -23, -38, 75, -39, -72, 47, -47, -54, 54, 29, -43, 33, -74, 36, -33, 21, -41, -50, -22, 57, -4, 48, 75, -25, 22, 45, -18, 48, -17, 11, -75, 33, 48, 73, 69, 49, 42, -55, 70, 21, 47, -51, -24, 46, 61, 18, -10, -56, 44, 43, 75, -38, 13, 72, 12, -43, 39, 67, -72, -54, 2, -74, 52, -26, 75, 46, -54, 41, 64, -62, -14, 35, -37, 36, 3, -54, -22, 68, -37, -54, 33, -40, -19, -32, -43, 69, 1, 71, 60, 4, -60, -15, 5, 67, 32, 2, 35, 53, -32, 21, 67, 27, -22, -46, -13, 57, -25, 41, 49, 11, 60, 5, 47, -36, 48, -72, -43, -27, 72, -61, 50, -66, -1, -22, 75, -44, 55, 32, -67, -53, -22, 75, 48, 29, -49, -41, 10, -1, 73, -18, -65, 56, 62, 57, -58, 32, 58, -26, -72, 52, -12, 53, 62, 61, -45, 59, -59, -67, 15, -53, -47, 66, -53, -75, 20, -29, -42, -46, 46, -47, 9, 54, -69, -7, 35, -52, -50, 15, -5, -47, -11, 57, -72, -27, 42, -43, -44, 56, -35, 47, -73, -9, 37, -53, -10, -21, -8, 21, 7, -38, 47, -60, -62, 54, 7, 46, 75, 30, -15, -7, 56, 47, -26, 59, -55, -62, -62, -24, 67, -22, -55, 67, 43, 56, -61, -43, -41, 4, 53, 41, 39, 24, 55, 52, 0, -14, 22, -2, -60, -71, 66, 71, 51, -38, 52, 71, -27, 66, -30, -36, -34, -10, -45, -67, -32, -33, -37, 3, 46, -62, -34, 9, 36, -55, -15, -42, 6, -69, 31, 19, -65, 19, 12, 60, 56, -11, 55, -47, -23, -51, -10, 18, 13, 21, 25, 56, 61, 63, -19, 32, -74, 23, -37, 37, 43, 22, 70, -28, 28, 24, 64, 37, -33, 1, 19, -54, 63, -2, -28, -36, 21, 38, 55, -42, -19, 4, -64, -36, -8, -7, 71, -9, -62, -43, -50, 54, 54, -58, -50, 4, 41, -63, -37, -69, 11, 57, -48, -4, -20, -3, 35, 74, -41, 12, -46, 13, -59, -35, 53, 8, 31, 46, 72, 42, -73, -54, 21, 54, -37, 44, -17, -71, 56, 19, -65, -9, 1, -40, 60, 54, 32, 19, 52, 65, -44, -70, 0, -30, -32, -23, 51, 73, -54, 47, 39, -54, 68, -16, -75, -45, -49, -19, -43, -69, 75, -35, -4, 0, 0, -20, -24, -45, 73, -48, -56, -49, -45, 17, -4, -3, 70, -29, -8, -62, -60, -45, -41, -68, 13, -43, -40, 39, 13, -9, 43, 11, 31, -39, -67, -46, 17, -15, -18, 12, 10, -1, 36, 39, -60, -44, -40, -68, 0, 25, -55, 13, 53, -20, 18, -12, 10, 51, -51, -52, -34, 68, 34, 71, -49, 42, -53, 41, -51, 4, -23, 35, -75, -63, -2, -60, -34, 31, -52, 39, -22, -34, -24, -45, 19, 69, 19, -46, 45, 43, -23, -67, 33, -67, -72, 60, 48, -52, 25, 73, 27, -75, 30, 25, -63, -50, 41, -23, 54, 62, -60, -44, -48, -8, -14, 47, -17, -73, -75, -50, 46, -25, -41, 1, -19, -40, -15, -47, -16, -67, -52, -67, -67, 51, 34, -57, -75, -3, -5, 54, -17, 9, -66, 8, -75, -6, -21, -19, -4, -23, 7, -36, 25, 39, 41, -70, 74, -52, -43, -18, -44, -22, -9, -38, -46, -53, -19, -48, 19, 51, -69, -74, -16, -62, 7, -18, 5, 62, 37, -74, -39, -34, -35, 62, -71, -72, 67, -75, -48, -54, -19, -17, 0, 45, 19, 29, 67, 75, 54, 10, 48, 58, 9, -45, 72, -62, 10, -1, 73, -31, 0, -41, 10, 39, -57, 12, 42, -68, 13, 69, -46, 69, -25, 29, 38, 69, -20, 27, 66, -42, -41, 38, -59, 41, 68, -65, 54, 1, 9, 52, 45, -66, -65, -20, 46, -47, 65, 12, -40, 2, 4, -11, -7, 54, -60, -47, 45, -5, 55, 35, 29, -64, -3);
    signal scenario_output : scenario_type :=(-21, 31, 61, 0, -88, 20, 48, -18, -5, 1, 54, -59, -75, 55, 0, -17, 18, 27, -30, 19, 49, -44, 1, 59, -51, -74, 77, 30, -19, 8, 9, -51, -64, 73, 35, -40, -17, -22, 51, 62, -18, -6, 24, -75, -63, 27, -2, 46, 34, -11, -24, -6, -37, -22, 32, 2, 14, -24, 57, -4, -12, 65, -60, -52, 3, 90, -5, -12, -22, -45, 71, -44, -51, 76, -26, -21, 80, -7, -64, 24, -22, 21, -2, -79, 111, 6, -52, 11, 4, 1, 3, 18, -65, 58, 52, -61, 58, -45, -51, 9, 20, 0, -53, 85, 49, -59, -26, 18, 43, 17, -69, -66, 39, 18, -31, 17, 26, 25, 27, -56, -62, 32, 47, -17, -18, -9, 55, 13, -54, 2, 26, -31, -21, 108, -62, -58, 46, 21, -41, -18, 41, -20, 6, 59, -4, -3, -12, -68, 41, -7, -30, 68, 24, -73, -38, 3, 27, -2, -1, 85, -1, -63, -39, 0, 20, -9, 30, 47, 13, 9, -63, -35, -12, 55, 2, -12, 49, -13, -55, -42, 89, 22, -83, 4, 61, -35, 9, -22, -17, 28, -51, -15, 56, 2, -37, 78, -9, 13, 36, -88, 23, 61, -32, 13, 3, -10, 21, -57, -23, 52, 11, -44, -35, 40, 47, 26, -85, -31, 4, -11, 90, -68, -3, 32, -70, 95, -23, -55, 109, -13, -7, 18, -42, -21, 29, -37, -29, 31, -5, 57, -27, -80, 13, 25, 71, -46, -57, 96, 9, -52, -2, -14, 11, -26, 0, 55, 41, 0, -91, 57, 5, -98, 57, 53, -5, -47, 40, -36, -17, 37, 0, 65, -45, -75, 2, 24, -35, 58, -11, 0, 5, -37, 98, -5, -43, 6, -41, 21, -20, -19, 59, -36, 20, -21, 41, 11, -70, 82, -25, -63, 3, -2, -18, 49, 11, -36, 76, -2, -70, -25, -4, 25, 51, -41, 42, 6, -35, 2, 7, 57, -20, -22, -66, 0, 45, 62, 9, -112, 34, 93, -66, -69, -18, 25, 71, -29, 13, 32, -10, -53, -13, 94, -28, -75, 77, 11, -69, 41, 12, -38, -12, -4, 27, 7, -5, -15, -15, 3, -17, -3, 76, 31, -96, 59, 56, -5, -61, -18, 28, 13, 39, -97, 21, 8, -62, 78, 0, 3, 4, -77, -32, 82, 5, -3, -17, 1, 91, -60, 27, -39, -39, 105, -34, 0, 49, -68, 13, -14, -87, 45, -21, 45, 39, -19, 55, -3, -30, -38, 21, -48, -23, 80, 11, 7, -37, 12, 28, -61, -21, 31, 8, -61, 26, -1, -62, 56, 21, 44, 18, -38, -24, 19, 4, 10, 23, -55, 34, -31, 19, 34, -79, 18, -1, -43, 4, 71, -31, -75, 12, 37, 48, -1, 0, -36, -2, 46, 17, -70, 2, 31, 0, -21, -55, 5, 79, 58, -49, 22, -66, -5, 31, -34, -6, 11, 32, -2, -25, 2, 31, -15, -46, -29, 95, 40, -68, 3, -1, -51, 23, 89, -17, -61, -44, 36, 29, 36, 5, -108, 60, 25, 0, -41, -4, 104, -34, -57, -10, 51, 55, -89, -74, 116, -10, -86, 47, 31, 8, 24, 3, -58, 24, -13, -31, 69, 22, -91, 14, 26, -86, 53, 32, 25, 8, -60, 39, -26, -8, 28, -83, 47, 25, -42, 32, 14, 4, -34, -42, 34, -32, 52, 65, -7, -52, -58, 83, -52, -34, 78, -47, 15, -5, 9, 38, 2, -27, -36, 2, -60, 82, 7, -8, -1, -11, 19, 10, -6, -12, -28, 4, 65, 22, -18, -30, -32, 34, 29, -82, 2, 82, 3, -95, -8, 9, 53, -28, -13, 21, -49, 38, 79, -19, -62, -12, -30, 45, 88, -34, -79, 81, -29, -12, 102, -53, -22, -40, -14, 96, -34, -9, 71, -32, 27, -76, 1, 80, -104, -9, 76, -19, -82, 44, 73, -57, 8, 66, -103, 7, 28, -72, 69, -2, -59, 37, 57, 4, -3, -46, 9, -18, -56, 57, 63, -51, -18, 68, 5, 12, -56, -6, -8, -28, 18, 44, 46, -85, 1, 56, 9, 29, -104, -10, 23, -51, 6, 61, 64, 1, -72, -37, 94, -19, -91, 46, 38, 2, 4, -43, 12, 57, -73, 6, 27, -56, 76, -59, -5, 54, -3, 28, -52, 27, -5, -25, -22, 0, 56, -69, 3, 71, 4, -13, -37, -64, 10, 91, 49, -96, -43, 83, -62, -2, 70, -32, -35, 9, 41, -42, -44, 39, 73, 12, -42, -17, -15, 42, -18, -69, -22, 72, 92, -15, -28, -61, 52, -19, -81, 103, -27, -9, 53, -70, 11, -10, 10, 63, 1, -58, 21, 65, -21, 5, -12, -44, -13, -27, -21, 58, -6, -41, 42, -7, -36, -10, 45, -5, -51, 79, 74, -57, -21, 12, 7, -35, 1, 39, -83, 5, 69, 49, -40, -41, 75, -56, -82, 41, 7, -10, 79, 0, -29, 9, -7, 41, -2, -51, -77, 81, 1, 0, 22, -21, 35, -85, -31, 14, 47, -25, 20, 26, -64, -21, 97, -11, -75, 14, 6, 43, 1, -1, -44, -29, 95, 57, -100, 6, 5, -64, 64, 8, -65, 90, -12, -29, 8, -68, 99, 31, -70, 9, 57, -25, -10, 43, -13, -91, 57, -6, -46, 60, -29, 20, 28, -20, -37, 62, -38, -30, 0, 5, 91, -68, 4, -11, -96, 103, 9, 4, 21, -39, 34, -34, -42, 23, -11, 30, 46, -87, 49, -2, -27, 18, 18, 2, -3, 5, -71, 72, 63, -71, -10, 39, -2, -27, 4, 34, -40, -72, 40, 69, 0, -36, -73, 69, 73, -82, 12, 3, -37, 38, 5, -63, 56, 21, -61, 55, 3, 1, 11, -22, -47, 2, -4, 38, 88, -110, -15, 43, -71, 25, -18, 42, 76, -92, 25, 34, -41, 12, 39, -56, -61, 46, -9, -25, 51, 38, 27, -35, -51, 41, 28, 11, -68, -63, 73, -5, -60, 36, 19, -17, 37, 24, -64, -1, 68, -65, 34, 26, -52, 78, -56, 23, -10, -42, -3, 38, 19, -89, 4, 56, 65, -76, -41, 107, -29, -77, -8, 22, 47, -11, 29, -27, 10, 74, -29, -32, 32, 3, -10, 3, -30, -42, 3, 49, 4, 2, -20, 22, 24, -19, -8, -23, 36, -51, -26, 7, -39, 56, 8, 8, 64, -53, -111, 99, -4, -27, 65, -82, 0, 32, 11, 58, -9, -72, 19, -6, 38, -2, -91, 64, 64, 11, -73, 13, -37, -9, 110, -76, -43, 27, -43, -1, 63, -42, -34, 64, 42, 4, 2, -48, -54, 37, -10, 26, 53, 9, -70, 2, 4, -53, 68, -38, -39, 83, 66, -76, -13, 62, -21, -59, -40, 48, 28, 4, 7, 12, -24, -42, 40, -43, 1, 78, -28, 11, 14, -64, 18, 58, -83, 25, 6, -39, 97, -31, -41, 48, 22, -60, 3, 4, -30, 72, -57, -89, 76, 39, 11, 52, -91, -34, 3, 22, 22, -22, 37, 35, -65, -58, 92, -37, -52, 77, 57, -68, -43, 32, -18, -38, 64, 72, -35, -53, 35, 15, -32, 0, -32, 2, 25, -8, -54, 31, 15, -31, 8, 51, 2, -58, 15, -38, 18, 52, 41, -37, 6, -5, -2, -10, -48, 85, -51, -58, 7, 75, 47, -22, -37, 39, -22, -11, 30, -77, 23, 22, 1, 32, -38, 27, -25, -42, 100, -10, -76, 26, 83, -72, -88, 82, 4, -20, 34, -44, 28, 40, -58, -10, 12, 13, 6, -5, 5, 11, 49, -85, -52, 52, 35, 25, -56, 31, 2, -69, 22, 35, -39, -26, 76, -17, -53, -28, 73, 68, -74, 14, -7, 2, -20, 8, 19, -15, 1, 24, 21, -83, 54, 56, -32, 0, -9, -66, 9, 82, -24, -78, 8, 46, 8, -46, 30, 63, -77, 17, 17, -15, 7, 9, -11, -11, 18, 7, -27, 17, 29, -7, -43, -26, 47, 32, -24, -94, 81, 72, -9, -53, 17, -2, -7, 25, -52, 46, -45, 7, 39, -29, 13, -64, -17, 92, 10, 0, 10, -109, 41, 19, -25, 87, -6, -68, 28, -35, -47, 90, 37, -35, -77, 54, 72, -87, -31, 44, -63, 35, 30, -21, 6, 24, 25, -12, 25, -54, 8, 10, -46, 27, 27, -49, 3, 22, -6, 10, -13, -31, -10, 23, 20, 23, -28, -17, 47, 27, 6, 6, -28, -54, 4, -24, -28, 6, 75, -23, -43, 83, -15, -69, 1, 14, -30, 96, 13, -13, 15, -90, -46, 95, 25, -25, 5, 15, -23, -61, 68, -20, -53, 19, 17, 43, -25, -12, 75, -62, -14, 27, 21, -29, -42, 24, -39, 62, -17, 1, 48, -24, 24, -1, -20, -38, -27, 75, 69, -53, -74, 25, 39, -37, 22, 77, -87, -91, 65, 75, -43, -60, -5, 90, -2, -46, 2, -19, 13, -13, -17, 40, 75, 4, -51, -32, -36, 31, 18, 36, -19, -55, 63, -4, 40, -27, -36, 64, -9, -80, 31, 57, -55, 26, 35, -34, -19, 37, -53, -6, 22, -72, 56, -14, -64, 95, 39, -98, 15, 79, -64, -2, 25, -5, 12, -44, -32, 90, -2, -40, 8, 27, 15, -46, 78, -63, -55, 36, 61, 1, -79, -23, 42, 66, -61, 1, 49, -22, 34, -45, -51, 80, 38, -25, -13, -60, 39, 63, -81, -49, 19, 38, -44, 34, 17, -99, 87, 46, -62, 40, 49, -31, 13, 1, -59, -25, 2, -31, 65, 13, -77, 37, -18, -14, -11, 58, 38, -82, 11, 66, -45, 35, -5, -70, 70, -11, -34, 21, 35, 34, -52, -5, 23, -37, -23, 55, 26, -43, 48, -20, -6, -29, -5, 90, -70, 8, 36, -36, 58, -63, -57, 31, -52, 29, 55, -2, 17, 42, -73, -39, 76, -12, -42, -32, 59, 42, -89, 0, 0, 47, 69, -5, -71, -27, 83, -29, -21, 7, -39, 13, 34, -6, 25, 3, -66, -9, 19, -52, 12, 38, 24, -43, 24, 93, -79, -2, 21, -36, -25, 22, 34, -71, 21, 51, 12, -8, -66, -6, 86, 4, -104, 31, -3, 34, 14, -70, 25, 13, -5, 13, 53, 17, -8, -12, 17, -68, -13, 19, -12, 46, 45, -90, -1, 62, -42, 38, -82, 26, 6, 3, 31, -95, 37, 28, -58, 27, 71, -32, -47, -27, 0, 5, -28, 83, 81, -9, -73, -23, 6, 21, 25, -79, 69, -1, -18, 53, -100, 36, 56, -91, 43, 63, -52, -31, -18, 23, -26, 31, 103, -76, -82, -8, 38, 0, -34, 9, 102, -19, -12, 18, -86, 7, 48, -39, 9, 34, -12, 44, -40, -68, 88, -23, -1, 37, -56, -18, 38, 29, 12, 26, -23, -70, 18, 15, -92, 97, 23, -81, -10, 8, 25, -5, -1, 76, -25, -81, 0, 73, 51, -63, 30, 25, -64, 29, 41, -9, 7, -9, -72, 45, -5, -7, 88, -98, -77, -4, 89, 37, -106, 79, 44, -59, -19, -46, 15, 44, -38, 19, 9, 10, 85, -73, -47, 17, 64, -8, -100, 77, 66, -62, 10, -27, -45, 76, -35, -32, 74, -55, 0, 99, -90, -43, 41, -19, 1, 38, 24, -14, -57, 54, 14, -82, -14, 52, 48, -82, 46, 57, -7, 24, -92, 2, 83, -27, -29, -62, 71, 18, -114, 75, 93, -72, -80, 26, 19, 7, 66, -65, 15, 4, -11, 35, -99, 86, 63, -25, -89, 20, 28, 13, 22, -63, 38, -8, -66, -15, 42, -13, -17, 38, 58, -32, -9, -24, -8, 9, -15, 57, -55, 0, 63, -65, 9, 100, -95, -11, 70, -73, -12, 103, -60, 8, 36, -20, 1, -29, -31, 22, 65, -53, -24, 13, 24, 53, -12, -74, -25, -27, 73, 6, -24, 26, -40, 7, -6, -21, 87, 40, -73, -17, 28, 2, -32, 68, -17, -31, 39, -54, 14, -28, 6, 77, -15, -56, 41, -26, -41, 103, -55, -53, -1, 29, 62, -60, 41, 52, -61, 38, -23, 0, -3, 6, 3, -37, 75, -17, -44, -20, 43, 57, -49, -37, 45, -70, 17, 64, -98, 2, 35, -41, 37, 11, 14, -17, -25, 56, 30, -66, -17, 10, 20, 88, -92, -64, 73, -41, 31, 6, -64, 103, -71, 20, 41, -44, 85, -55, -66, -12, 36, 56, -49, -38, 90, -37, -54, 63, 17, -22, -2, -1, -13, 42, -45, 6, 68, 4, -9, -13, 31, -52, -48, 98, -56, -6, 75, -85, -37, -13, -3, 90, 20, -32, -39, -1, 38, 14, -48, -30, -8, 38, 57, -18, -30, 29, 8, -78, 59, -25, 23, 69, -79, -1, 31, 0, -8, -25, 31, 39, -39, -61, 39, -19, -4, 90, -21, -53, -6, 41, 3, -13, -10, -28, -34, 69, -18, -46, 106, 17, -51, 38, -25, 2, 32, -107, 28, 0, -19, 39, 41, -59, -20, 81, -83, 0, 38, 6, 34, 30, -40, -52, 15, 39, 7, -17, -4, 8, -43, -7, 26, 15, 7, -1, 43, -94, 26, 49, -91, 6, 88, -47, -53, 70, 7, -3, -44, -44, 25, -9, -35, 76, 27, -19, 24, -56, -12, 0, 44, 31, -8, -17, -45, 18, -18, -22, 40, -12, 5, 61, -4, -15, 31, -39, -58, 42, 48, -11, 0, -36, -24, 75, 40, -87, -34, 65, -54, 40, 66, -99, -18, 57, -27, 29, 54, -23, -82, -18, 74, 31, -69, -20, 38, -58, 32, 69, -15, -8, -34, -15, 44, 54, -55, -5, -11, -89, 40, 22, 64, -25, -51, 45, 26, -56, -36, 82, 6, -7, -44, -6, 20, -1, -46, 40, 49, -17, 20, -54, -24, 72, 41, -92, 38, 6, -99, 5, 9, 30, 30, -36, 24, -20, 8, 52, -78, -2, 2, 42, 75, -44, -51, -13, 63, 9, -86, 28, -7, 22, 64, -32, 8, -8, 6, 24, 0, -93, 28, 9, -61, 61, -24, -36, 40, -14, -5, 76, -43, 17, 25, -56, -24, 60, 41, -69, -40, 65, 46, -47, 0, 20, -61, 6, 11, -55, 31, -9, -31, 43, -21, 18, 83, -46, 5, 9, -41, 21, -51, 52, 14, -22, -4, -8, 39, 13, 34, -3, -7, -10, -30, -8, -13, 21, -20, -22, 80, -11, -11, -41, -78, 79, 64, 2, -55, -18, 9, 13, -19, -38, 64, -4, -61, 62, -11, -25, 97, -92, -3, 63, 7, -34, -56, 18, -35, 14, 85, 46, -86, -17, 1, -53, 40, 70, -49, -13, 51, -41, 1, 6, 54, -45, -86, 13, -6, -5, 81, 70, -76, -15, 44, -66, 40, 78, -48, -83, 3, 34, 51, 28, -91, -57, 87, 38, 12, -54, -66, 64, -8, 48, -38, -42, 3, -35, 62, -23, -14, 30, 42, 41, -95, -23, 82, 54, -57, -54, -28, 32, 93, -90, -46, 111, -37, -70, 61, -24, -34, 87, 19, -20, 21, 2, -62, 2, 81, -23, 0, -26, -83, 63, -8, -63, 17, 74, -9, -40, 19, -38, -3, 89, -15, -48, 92, -56, 13, 14, -58, -1, -10, -14, -22, -9, 79, 4, -5, 49, 2, 13, -92, -56, 55, -7, -27, 53, 66, -18, -75, -26, 52, 31, -70, 60, -20, 17, 26, -117, 36, 58, -26, 4, 44, -51, 18, 10, -25, 30, -54, 1, 23, -53, 37, 57, -62, 29, 21, -88, 9, 34, -21, 43, 68, -70, -9, 70, -52, -5, 63, -19, -35, -53, -14, 99, -13, 3, -3, -17, 34, -59, -12, 36, -2, 24, -14, -42, 53, -17, -13, 41, 17, -15, -4, -28, 45, -17, -71, 15, -23, -27, 90, 28, -79, -11, 12, 37, -29, 11, 22, -17, 63, 7, -70, -26, 30, 1, 44, -49, 10, 27, -11, 49, -100, 6, -3, 36, 79, -71, -56, 53, 32, -79, -27, 64, -3, -12, -7, -10, -1, -9, 107, -51, -91, 37, 10, 28, 43, -56, 0, 52, -30, 9, -34, 5, -5, -35, 44, 52, 4, -15, 18, -74, 18, 78, -9, -73, -46, 94, 3, -46, -4, 0, 13, -6, 15, 47, -68, -53, 103, 18, 0, -14, -62, -11, -32, 23, 42, 8, -12, -41, -6, 92, -1, -102, 82, -12, -61, 17, 58, 54, -29, -36, -36, -14, 42, 93, -103, -2, 61, -114, 40, 40, -39, 69, 5, -49, 3, -40, -42, 78, 7, -46, 61, 1, -12, 12, -10, 34, 26, -41, 0, -5, 35, -60, -22, 104, -103, 9, 77, -62, 34, -18, -1, 14, -58, 6, 52, 31, -34, -75, 0, 80, -13, -47, -5, -26, 49, 95, -104, -9, 52, 4, -12, -48, 78, -35, -78, 110, -27, -110, 48, 93, -14, -60, 0, 32, 54, -60, -19, 17, -26, -15, -35, 74, 23, -61, 71, -15, -78, 79, 61, -24, -7, -45, -49, 51, 7, -14, 30, -18, 5, -32, -34, 102, -5, -37, 48, -65, 38, 3, -47, 13, -32, 32, 65, -9, -7, 22, -5, -64, -8, 54, 21, -37, 9, -5, -99, 20, 69, 18, 4, -37, 6, -9, -47, 2, 43, 92, -63, -6, -17, 22, -17, -49, 78, -64, -36, 47, 49, 45, -15, -47, 10, 1, 25, 1, -23, 37, 18, -42, -31, 18, 30, -46, 9, -14, -45, 77, -61, 26, 47, -75, 51, 4, 8, -7, -31, -28, 35, 40, -93, 20, 77, 31, -89, 11, 52, -113, 53, 45, -46, 23, -43, -17, 88, -54, -29, 41, 0, 43, -46, -41, -8, -20, 78, -20, -26, 43, -49, 10, 59, -7, -81, 47, 19, -59, 41, 49, -39, -15, -11, 25, 92, -55, -77, 69, 0, 1, 0, -88, 43, 41, -38, 11, 46, -74, 13, 19, -52, 76, 25, -80, -42, 57, 56, -45, 21, -14, 27, -19, -31, 13, 4, 62, -42, -48, -3, 71, 42, -26, 4, -4, -75, -10, -13, 62, 6, -19, 80, -26, -31, -4, 2, 35, -59, -27, -8, 49, 69, -94, -57, 37, 6, 62, -35, -13, 13, -39, 76, -57, -39, 59, 28, -24, 25, 36, -52, -58, 38, 1, 28, -13, 0, 31, 20, -59, 2, 10, -7, 71, -86, -61, 87, 34, -24, 77, -93, 8, 36, -14, -51, -4, 44, -23, -4, -40, 12, 28, -5, 30, 54, -70, -74, 52, 73, -76, -2, 74, -69, 13, 11, -41, 62, -36, 13, 58, -71, -56, 43, 57, 19, -5, -38, -24, -28, 45, 24, -12, -36, 38, 37, -96, -28, 54, 48, 21, 0, -43, -17, 64, -54, -3, 20, 5, -17, -77, 66, -1, -21, 0, -31, -2, 83, 19, -26, -36, -22, -2, 36, 49, -73, -32, 66, -14, 18, 27, -83, 17, 72, 11, -53, 41, 5, -30, 47, -11, -83, -20, 100, -15, -41, 69, 1, -48, 0, -27, 3, 66, -27, -47, 5, 10, 7, 51, 15, -62, -32, 42, 64, -74, -35, 32, -32, -29, 3, -4, 47, 8, -23, 38, 11, -45, -4, 11, 15, -25, -11, 21, 18, 72, -27, -66, -10, 0, -13, -11, 27, 41, 30, -19, -7, -3, -8, 71, -56, -2, 62, 11, -86, -49, 51, 14, -3, 23, 51, -77, -90, 39, 28, 39, 0, -86, -27, 80, 5, -61, 70, 30, 0, 9, -80, 12, -19, 25, 63, -76, 45, 14, -60, 47, 53, -9, -25, -39, 37, 0, -28, 59, -73, -86, 97, 14, -80, 73, -17, -52, 10, 49, 0, -102, 61, 9, 2, 42, -52, -46, 79, 80, -32, -70, 37, 40, -83, 9, 1, -43, -9, 87, -7, -80, 3, 68, 47, -77, 31, 30, -22, 41, -27, -21, 53, 8, 8, -37, -36, -45, 25, 43, -74, -8, 83, -55, 11, 112, -47, -73, -44, 74, -8, -72, 106, -7, -93, 43, 24, 46, -38, -85, 89, 20, 3, 30, -60, 37, -28, 12, -7, -114, 59, 4, -9, 9, -28, 25, -12, 37, 41, -57, 2, 30, 2, -23, 26, 18, 14, -36, -43, 87, -11, -65, 14, 12, -35, -42, 26, 46, -46, 0, 45, -7, 6, 36, -2, 0, -49, 6, 35, -8, -52, 39, 22, -51, 38, -66, -5, 30, -13, 63, -15, -1, -4, 0, 12, -63, 74, 17, -15, 46, -75, -59, 35, 41, -43, 35, 42, -93, 42, 57, 10, -11, 5, -58, -40, 19, -34, 45, 30, -23, -4, 36, -27, -8, 37, -18, -49, 0, -2, 46, 24, -74, -10, 37, 79, -57, -13, 8, -18, 24, -46, 15, 12, -62, 47, 66, -63, 38, -1, -11, 13, -5, 22, -17, 8, -48, -34, 46, 38, -31, -12, 63, 1, -25, 9, -10, -58, -27, 88, 12, -1, -44, -82, 124, -20, -31, 77, -63, 4, 74, -53, -94, 71, 57, 2, -56, 30, -31, -7, 70, -69, 1, 18, -45, -23, 8, 35, 5, -15, 12, 41, -18, -56, 96, -30, -53, 62, 22, 17, -45, 8, -38, -26, 57, 21, -24, 1, 49, -59, 21, -15, 6, -1, 3, -36, -24, 13, -21, 93, -4, -95, 22, 86, -41, 4, -34, -71, 43, 99, -54, -112, 110, -5, -28, 57, -74, -29, 36, 64, 22, -53, -37, 27, 55, -55, -6, 29, -42, -3, -9, 62, 8, -97, 41, 79, -3, -14, 28, -47, -27, 82, -49, -26, -31, 34, 117, -108, -82, 42, 70, 25, -11, -55, -36, 43, -21, 48, 52, -42, -46, -47, 20, 51, -34, -48, 20, 74, 44, -63, -62, 40, -5, 0, -9, -32, 36, 82, -27, -46, 36, -52, 0, 1, -14, 58, 22, -14, 13, -12, -58, 57, 29, -35, -3, -2, 25, 12, -18, -18, -51, 28, 0, -54, 31, -31, 24, 70, -61, 17, 22, -48, 80, 0, -24, -25, -32, -1, 47, 72, -12, -99, 37, 13, -22, 11, 9, 25, -83, -5, 94, -22, -107, 97, 35, -96, 66, 60, -28, 23, -14, -95, 0, 39, 17, -43, -5, 95, -47, -44, 53, 47, -35, -19, -25, -58, 85, 74, -32, -90, -21, 63, -24, -13, 27, 10, 20, -19, -17, 10, 6, -53, 5, 93, -9, -89, 69, 3, -107, 24, 46, 58, -38, -75, 39, 22, -22, 12, -12, 58, 9, -31, 9, 4, -26, -74, 18, 82, -3, 1, -13, 1, 58, -10, 5, -43, -77, 53, 48, -73, -32, 8, -13, 17, 25, 3, 41, 3, 36, -63, -27, 43, 14, -17, -63, -8, -1, 44, 52, 17, -43, -54, 39, 9, -61, 25, 54, -27, -29, -4, 10, 25, -13, -1, 39, 30, -89, -7, 36, 34, 41, -104, -10, 56, -31, 18, 24, -11, -26, -11, 5, 17, 24, 24, 28, -15, -40, -5, -45, 18, 80, -35, -45, -26, -14, -25, 98, -14, -32, 43, -72, 9, 29, 7, 43, 19, -64, -20, 9, -3, 56, 15, -77, -9, 60, -49, -23, 0, 35, 18, 21, 3, 7, -22, -45, 105, -51, -35, -23, 28, 97, -96, -51, 13, 24, 80, 11, -15, -30, -70, 1, 1, 38, 14, -5, -9, -36, 81, -34, 22, 8, -105, 46, -6, -14, 1, -34, 48, 53, -58, -8, 38, -42, 27, 29, 5, 17, -46, -10, 74, -27, -6, -34, 30, 5, -38, 20, -29, 42, -13, -7, 31, -4, 14, 26, -18, 14, 10, -58, -41, 64, 20, -25, 45, -44, -86, 54, 58, -21, -66, 24, 62, 12, -9, 4, -71, -49, 115, -11, -3, -10, 1, 25, -17, 40, -63, -11, 56, -76, 40, 13, -121, 62, 99, -97, 21, 11, -44, 85, -32, 21, -5, -60, 56, -13, -77, 73, 48, -75, -25, 43, 22, -24, -44, 31, -8, 6, 0, 25, 63, -72, -68, 55, 78, 7, -18, 7, -70, -40, 66, 9, -19, -53, -26, 15, 23, 7, -21, -37, 44, 41, 9, -41, 14, 72, -9, -78, -34, 98, 58, -82, -64, 8, -28, 17, -5, 64, 3, -72, 26, 46, 51, -14, 17, -68, -89, 40, 28, -17, -15, 77, 19, 11, -54, -54, 85, 20, -20, -60, 30, 34, -30, -53, 21, 54, -59, 40, 7, -56, 78, 32, -99, 37, 41, -104, 61, 40, -62, -18, 21, 54, -54, -46, 64, -20, 11, 37, -88, -8, 65, 34, 26, -77, 3, 45, -25, -30, -46, 93, 22, -77, 12, 54, -40, -79, 88, -3, -36, 26, -21, -13, 57, 36, -59, 9, 35, -25, -87, 62, 51, -21, 9, -37, 35, -10, 10, 8, -42, -12, -8, -19, -2, 98, 12, -21, -70, -11, 88, -19, 14, -45, -8, 70, -10, -46, -31, 27, 11, -5, -19, -23, -27, 79, 28, 7, -19, -49, 18, 24, 26, -12, 27, -66, -3, 40, 0, 37, -83, 0, 19, 19, 65, -102, 1, 52, -37, -25, -52, 87, 54, -69, -48, 49, 8, -20, 57, -14, -48, -34, 11, 64, 66, -72, -90, 61, 57, 21, -35, 0, 18, -18, 40, -28, -96, 43, 2, -44, 106, -48, -42, 49, -9, 20, -35, 20, 19, -88, 6, 60, -32, 19, 38, -79, 60, 35, -18, 25, -32, -32, 23, -13, -49, 43, 46, -30, -43, 47, 57, -73, 24, 9, -23, 14, 27, -37, -76, 51, -36, 21, 89, -46, -46, 11, 6, -12, 48, -10, 13, 14, -43, 40, -23, 39, -29, -63, 2, 37, -11, -72, 77, 98, -61, -36, 25, -32, 14, 40, -6, 2, -25, -31, 68, 14, -17, -37, 25, 29, -47, 40, 42, -72, -32, 43, -55, 28, 69, -49, -42, 55, 8, -78, 43, 56, -3, -41, -65, 32, -26, 41, 12, -51, 30, -32, -10, -10, 45, -9, 18, 19, -81, 63, 32, 0, -25, 0, 47, -69, -26, 3, -34, 74, 14, 9, 41, -79, -32, 64, 42, -57, -1, 54, 20, -81, -86, 119, -7, -37, 1, 10, 89, -80, -12, 32, -86, 71, 12, -35, 2, -35, 81, -35, -51, 7, -26, 80, 17, -58, 60, -55, 15, 32, 4, 37, -53, -58, 22, 55, -8, 23, -21, -12, -36, -57, 111, -8, -95, 12, 69, -4, -21, 41, -38, 38, 23, -40, 7, 40, 31, -47, -100, 47, 71, 14, -28, -70, -20, -28, 79, 58, -4, -29, -68, 70, 23, -68, -48, 40, 35, -2, 57, -78, -48, 17, 48, 65, -21, -32, 14, 9, 6, 25, -55, -8, 41, 7, 11, -2, 0, 0, -34, 18, -56, 10, 66, -29, -55, 17, 9, -22, 39, -65, 12, 77, -48, -27, 52, -48, -61, 44, 73, -55, -40, 19, 44, 1, -85, 78, -1, -80, 57, 54, 27, 3, -23, 4, -29, 30, -1, -19, 31, -74, -61, 21, 95, -19, -2, 35, -48, -45, -32, 26, -11, 19, 26, 37, 19, -36, 3, 12, 12, -51, -19, 38, 60, -44, -68, 57, -37, 44, 13, -3, -28, -46, 20, 41, 69, -95, -10, 18, -49, 47, 22, -35, -46, 72, -2, -28, 35, 0, 8, -85, 63, 76, -44, 11, 51, -94, -41, 14, 37, 86, -100, -79, 40, 8, 75, -26, -60, 64, -32, 24, -21, -6, 97, -72, -20, -15, 10, 102, -18, -68, -71, 43, 93, -3, -53, 34, 11, 15, -61, -38, 100, -73, -1, 4, -39, 74, -48, 35, 4, -55, 57, -20, -39, 20, 22, 27, 5, -56, 39, -11, -36, 58, 31, -31, -37, -1, 0, -22, -6, 26, 55, -40, -21, 51, -39, -36, -9, 49, -25, -3, -4, 8, 87, -45, -57, 20, -18, 35, 53, 21, -64, -73, 79, 55, 5, -70, -32, 6, -3, 48, 35, -38, -82, 13, 103, -29, -19, -17, 17, 65, -22, -77, -14, 62, -32, 19, 61, -28, -36, 23, -10, 9, -47, -39, 65, 44, 1, -80, -34, -2, 59, 91, -62, 0, 12, -51, -7, -31, 46, -12, 32, 23, -90, 21, 63, 10, -72, 36, -21, 3, 38, -27, 14, -36, 66, -32, -76, 68, -22, -21, 42, 59, -23, -108, 61, 76, -44, -79, 46, 112, -94, -6, 21, -53, 12, -46, 75, 30, -34, 76, -56, -85, 48, 44, -5, -17, 11, 49, -87, 14, 26, -42, 75, -21, -14, 19, -31, -60, 48, 15, -83, 93, -15, -60, 44, -26, 28, -19, 26, 15, -55, -25, 19, 80, 19, -75, -27, 55, -48, 0, 46, -22, -18, -11, 68, 77, -103, -52, 15, 35, 54, -62, 18, 35, 6, -52, -77, 37, 17, 40, 34, -39, 34, -36, -46, 53, -24, 38, -27, -47, 39, -3, 44, -2, 5, 22, -40, 37, -52, -22, 72, 0, -63, -22, 36, 35, 13, -39, -37, 52, -1, -4, 37, -80, -40, 80, 61, -62, 10, 31, 21, -65, -58, 63, 41, -53, -25, 26, -40, 34, 4, -80, 35, 31, -11, 72, -23, -87, 28, 48, -55, 29, 43, -15, -48, 3, 61, 9, -35, -42, 65, -38, 5, 6, -82, 47, 40, 6, -59, 24, 39, -77, 59, 52, -24, -43, 10, 62, -19, -69, -1, 55, -39, -65, 39, -3, 49, -8, -81, 13, 39, 74, -24, -43, -29, 4, 91, 10, -78, -57, 35, 48, -22, -15, -8, 61, 51, -108, 35, 27, -66, 38, -46, 4, 61, -27, 25, 0, -37, 55, 11, -90, 39, -9, -43, 97, -5, -39, -5, 27, -6, 30, -34, -7, 11, -43, 56, 38, -18, -20, -22, -64, -3, 22, 31, 36, 13, -32, -54, 0, 0, 47, 3, 18, 37, -20, 21, -59, -35, -6, 57, 69, -88, -62, 60, 10, 5, 5, -40, 9, -38, 28, 37, -62, 54, 68, -5, -22, -56, -60, 65, 34, -10, -21, -40, 46, -40, -37, 79, 11, -44, 49, -30, -21, 76, 7, 11, -7, -77, -28, 92, -25, 2, 15, -66, 76, -30, -47, 30, 3, 6, -38, 62, -6, -60, 24, 15, 10, -13, -13, 22, 74, -100, 15, 51, -24, 45, -48, -31, 55, 35, -54, -58, 37, 49, -11, 1, -69, -37, 8, 26, 57, -27, -18, 48, 22, 3, -24, -55, -11, 70, -31, -71, 106, -41, -15, 79, 1, -43, -65, 81, -35, -3, 2, 4, 46, -9, 4, -22, -47, 13, 4, 8, -11, -13, 58, 6, 11, -80, -25, -21, 80, 31, -89, 75, 10, -86, 42, 14, -40, 89, -37, -48, 82, -40, -21, 14, -27, -14, -28, 17, 89, -22, -82, 77, 73, -27, -5, -27, 27, -54, -46, 110, -48, 1, 48, -14, -64, -20, 0, 6, 46, -40, -18, -3, 35, 48, -8, 9, 31, -15, -61, 7, 71, -35, -26, 54, -43, -32, 27, -39, 21, -13, -60, 109, -38, -8, 93, -103, -24, 68, 17, 0, 28, 19, -94, -25, 64, 5, -13, -10, -11, 31, -1, -54, 18, -28, -19, 69, 25, 7, -57, -62, 103, -6, -89, 89, -14, -18, 98, -42, -37, 22, -21, -8, 18, -4, -32, -25, 3, 41, 53, -9, -15, -38, -64, 94, 21, -82, 48, 70, -76, -7, 7, 3, 97, -81, 2, -8, -75, 78, 37, -2, -11, -73, 11, -17, 12, 72, -64, 38, 19, -102, 29, 94, -51, -32, 76, -29, 15, 9, -49, -38, -18, 48, 78, -56, -6, 79, -69, -61, 43, -9, -62, 12, 8, 39, -26, 47, -4, -69, 86, -7, -34, 1, -23, 23, 77, -56, -93, 92, 43, -51, 31, 44, -90, -1, 119, -99, -30, 48, -47, -7, 20, 2, -17, 31, 39, -21, -32, 32, 40, -61, -61, 7, 28, 3, 34, -2, -54, 74, -47, 12, 22, -14, 58, -69, 7, 40, -31, -45, 71, 30, -55, -17, 32, 36, 12, -17, -75, 0, 13, -53, 29, 44, -64, 60, 46, -7, -56, 12, 64, -103, 27, 62, 14, -28, -96, 45, -8, -39, 110, -49, -93, 56, 18, 49, -17, -53, 31, -3, 38, 23, -34, -19, -44, 31, 17, 5, 23, -40, 43, -49, -7, 46, 14, 8, 15, -58, -59, 5, 14, 31, -63, 35, 61, -18, -26, 44, 38, 0, -48, -11, 24, 27, -55, -17, 61, -41, 9, -28, -59, 30, 12, 21, 79, -60, -60, 95, -31, -3, -30, 6, 22, -93, 45, 62, -1, 14, 18, -54, 37, -34, -66, 64, -28, -8, 24, 31, -26, -75, 5, 2, 46, -2, 51, 9, -42, 11, -30, 63, -15, -59, 73, -19, -20, 4, -46, 2, 0, 60, 60, -76, -61, -5, 79, 0, -15, 17, -79, 69, 28, -71, -37, 71, 59, -102, -3, 17, -2, 80, -54, 2, 40, -93, 9, -1, 1, 54, -21, 22, 23, -51, -52, 53, 31, 24, -37, -72, 42, -4, -25, 51, 36, -64, 37, -18, -32, 9, -22, 102, -45, -53, 104, -29, -9, -22, -6, -6, 9, 82, 13, -56, -60, -17, -27, 63, 99, -64, -95, 30, 38, -8, -51, 78, 36, -13, -48, 2, 106, -73, -4, 57, 6, -13, -61, -1, 53, 20, -9, -28, 12, 25, -87, -68, 102, -25, -1, 93, -93, 35, -13, -28, 23, -63, 48, 59, -77, -1, 61, 25, -52, -56, 105, -46, -68, 20, 62, -15, -66, 52, 62, -51, -53, 88, -9, -64, -26, 10, 3, -5, 26, -28, 77, 25, -69, 37, -29, -12, 10, 36, 10, -43, 4, -19, 24, 23, 5, -22, 2, 71, -82, -20, 14, -24, 49, -13, 24, 0, 0, 27, 10, -65, -91, 89, 47, -46, -5, 22, 49, 2, -31, -31, -15, -47, 40, 96, -25, -43, -15, 0, 0, 14, -39, 15, -8, 7, 2, 14, 4, 1, 65, -94, -61, 64, 86, -13, -72, -12, 26, -24, -6, -23, 34, 64, -73, -11, 51, 13, 29, 32, -75, -58, 48, -26, 49, 17, 4, -37, -58, 29, -35, -11, 25, -8, 54, 0, -22, 93, -13, -82, -43, 89, -19, -5, 40, -70, -17, 68, 77, -102, 11, 2, -47, 38, -20, 2, 55, -17, -31, -1, -10, 45, -36, 17, 58, -96, 39, 56, -115, 25, 59, -43, -18, 64, -49, 2, 106, -69, -18, 70, -37, -30, 72, -61, -104, 52, 30, 40, 35, -91, -49, 23, 42, 3, 44, -10, -70, 81, 18, -51, -2, -29, 17, 66, 9, -8, -20, 24, -59, -40, 71, 15, -66, 11, 64, -62, -46, 7, -20, 77, 5, -66, -6, 43, 68, -76, -57, 19, -14, 53, 60, -39, 42, -13, -62, 74, -26, -82, 80, 1, -10, 41, -71, -56, 29, 83, -26, -35, 92, -27, -46, -14, 17, 35, 30, -28, -17, -25, -30, 78, 23, -59, -52, 69, 11, -1, 12, -14, 46, -21, -100, 58, -3, -81, 94, 4, 24, -24, -119, 115, 35, -53, -10, -37, 3, -2, 24, 75, -27, -93, 40, 107, -64, -7, 63, -32, 11, -37, -24, 36, 28, -9, -35, 25, 38, -55, -55, 63, 6, -61, 46, 41, 18, -77, -83, 21, 7, 34, 78, -20, -39, 29, -27, 27, 20, -76, 18, 6, 0, -27, 45, 31, -39, 30, -56, 1, 63, 1, -43, -41, 72, 0, -111, 93, 11, -103, 96, 19, -45, 58, 18, -63, -26, 11, -35, -27, 28, 72, -18, -80, 68, 22, -49, 29, 30, 28, -81, 5, 28, -37, 79, -31, -14, -9, -75, 110, -1, -90, 18, 85, -36, -73, 23, 26, 31, -29, -1, 82, -72, 0, -1, -2, 24, -53, 27, 55, -25, -53, 62, 0, -66, 6, 80, 6, 0, -83, 4, 108, -64, -88, 83, 8, -49, -22, 36, 90, -56, -49, 60, 4, -74, 59, 1, -48, 6, 28, 6, -20, -2, -41, -18, 19, 56, 61, -61, -58, 89, 53, -63, -65, -12, -1, 35, 25, -25, -11, 6, 26, 45, -46, -56, -5, -7, 37, 34, 2, -45, 62, -20, -49, 24, -60, 80, 77, -90, -71, 39, -1, -38, 66, 26, -72, 68, 61, -26, -49, -41, -20, 69, 92, -63, -98, 87, 38, -61, 11, 36, 25, -60, 39, -26, -38, 0, -57, 40, 0, -37, 60, 0, -52, 14, 22, 7, -27, -26, 93, 11, -90, 96, -12, -87, 30, 0, -18, 48, 48, -8, -4, -15, -45, 11, 47, 6, -8, 15, -63, -8, 90, -27, -5, 36, 7, -72, -68, 87, 10, -86, -10, 55, -12, -42, 83, -4, -43, 82, -47, -81, 74, 37, -7, 25, -38, -49, 30, 65, -58, -32, 57, 30, -37, -60, 68, 58, -42, 1, 34, -8, -86, 23, 46, -102, 4, -5, 9, 52, 57, -39, -10, 41, -93, 2, 45, -39, 39, 78, -86, 4, 43, -27, 35, 2, -68, -8, 62, 0, -7, -10, -9, 15, -7, 15, 27, -4, -78, -54, 69, -44, 21, 36, -22, 39, 36, -66, -91, 98, -12, -62, 79, 29, -69, 2, 34, -26, -5, -15, -1, -34, 61, 79, -15, -35, 2, 35, -63, 39, -41, -17, 109, -21, -70, -5, 40, -56, 18, 40, 21, 6, -2, 10, -54, -48, -8, 70, 15, -10, -55, 12, 61, 4, 4, -46, -10, 7, -34, 38, 25, -76, 44, 20, -73, -47, 104, 58, -103, 34, 5, -62, 40, -14, 40, 75, -62, -55, 30, 63, 20, -23, -10, -8, 0, -10, -52, -28, 87, 24, -100, 2, 60, 35, 0, -12, 8, 12, -46, -74, 24, 52, -42, 42, 58, -95, 27, -6, -40, 60, -55, 4, 11, 43, -4, -97, 36, 30, -11, -8, 56, -1, -8, 27, -57, 10, 12, -47, 4, 57, -30, 32, -2, -53, 77, 31, -14, -10, -64, -34, 25, -28, 61, 38, -72, -55, 51, 54, -42, 40, 61, -78, -49, 53, 36, 2, -44, -58, 68, 46, -2, -53, -6, -7, 1, 69, -89, 11, 35, -41, -40, 42, 42, 19, -28, -30, 74, 21, -65, -61, 82, -26, -23, 9, 24, 34, -97, -18, 82, -30, -78, 83, 3, 4, 76, -85, -15, -14, 39, 0, -75, 111, 17, -8, 40, -106, -17, 90, 25, -82, -79, 112, -22, 6, 9, -83, 41, -1, 10, -5, -28, 44, 52, -2, -40, 11, 47, -80, 0, 87, -82, -49, 61, 68, -60, -34, 98, -80, -53, 127, -76, -19, 105, -77, 10, -20, -24, 26, -18, -9, -3, 62, 31, -41, -30, 11, -26, -6, 43, -24, -53, 75, 11, 9, 30, -27, 0, -7, 25, -53, -14, 82, -74, -17, 8, 24, 51, -15, -36, -79, 83, 47, -14, 27, -85, -25, 17, -18, 58, 41, -43, 27, 2, -12, 58, -79, -15, 30, 26, -12, -20, 37, -66, 41, -5, -57, 66, 43, -51, -82, -12, 11, 56, 85, -96, -2, 57, -79, 0, 4, -38, 65, 9, -34, 78, -70, 22, 37, -35, 49, 21, -34, -25, -19, -17, 58, 35, -62, 15, -15, -56, 93, -5, -87, 64, 30, -92, -9, 68, -2, -26, 53, -52, 5, 19, 3, 68, -73, -45, 52, -26, -21, -1, 38, 46, -15, 6, -8, -56, 0, 64, 0, -17, -52, 46, 23, -17, -46, 13, 52, -52, 9, -30, 34, -10, -11, 63, -79, 51, -7, -22, 22, -32, -1, -49, 18, 70, 46, 8, -77, -42, 71, 35, -82, 20, 81, -59, 4, 31, -22, -56, -17, 74, 23, -94, -22, 10, 57, 13, -74, 73, -11, -51, 43, -36, 10, 58, -56, -30, 69, -45, 38, 6, -10, 89, -86, -19, 49, -85, 14, 8, -48, 89, 62, -24, 15, -53, -104, 72, 47, -61, 12, 36, 0, 34, 21, -80, -17, 75, -3, -61, -57, 36, 31, 45, -8, -28, 26, 15, 20, -73, -64, -5, -4, 87, 80, -99, -75, 90, 60, -28, -62, -14, 5, 45, 19, -81, -32, 91, 83, -31, -83, 47, -1, -26, -15, -9, 54, -13, 32, -58, 28, 53, -63, -64, 48, 18, -75, 86, -27, 10, 56, -91, -4, 61, -41, -8, 91, -75, -4, 62, 0, 22, 0, -88, -5, 68, 13, -62, -31, 43, -11, 0, -35, 38, 24, -5, 55, -29, -31, 47, 1, -89, -40, 86, 59, -80, -7, 37, -25, -13, -12, -1, -13, 78, 0, -20, 59, -99, 52, 1, -54, 42, -23, 46, -56, 26, 37, -1, 20, -111, 72, -2, -87, 10, 63, 86, -73, -30, 10, 10, 42, -24, 34, -62, -37, 32, 27, 0, -64, 80, -22, 19, -13, -20, 62, -73, 28, -12, -48, 23, -9, 1, 0, 14, 10, -22, -10, 48, 32, 0, -26, -15, -2, -15, 11, 49, 17, -48, -41, -26, 4, 52, -29, -5, 34, 7, 59, -74, 19, 6, -52, 11, -11, 63, 0, 21, -73, 14, 68, -43, 37, -73, -35, 10, 0, 90, -48, -72, 39, 1, -5, 24, 51, -14, -72, -5, -5, 76, 29, -98, -24, 92, 0, -37, 43, 23, -15, -32, 59, -61, -49, 74, -43, 4, 64, -18, -19, 14, 21, -2, 37, -75, -66, 88, -1, -45, 60, 13, -60, -20, 25, 25, -62, 49, -13, -19, 73, -31, -25, -1, 17, 34, -61, -1, 38, 3, -20, 18, 41, -113, 39, 53, -77, -24, 10, 32, 37, -37, -61, 89, 29, -34, 2, -10, 12, -11, -4, -47, 69, 54, -46, 0, -25, 27, -27, 13, 29, -46, 35, 45, -26, -38, -7, 7, 22, 2, -45, -51, 73, 2, -72, -7, 81, 18, -14, -17, 25, -23, -63, 96, 29, -91, -15, 7, 24, 45, 21, -32, -93, 77, -10, -5, 15, -17, 2, 39, -15, -41, -9, 36, 72, -85, -57, 41, 45, 13, 24, -39, 10, -19, -54, 42, -19, 20, 27, 28, -24, -41, -8, -6, 13, -17, -9, 9, 77, -9, -38, -48, 59, 39, -10, 19, -24, -48, -51, 25, 55, 63, -14, -24, -47, -46, -3, 24, 62, 24, -36, -53, -15, 46, 31, -22, 31, 21, 5, 15, -78, -35, 79, -41, 7, 66, -21, -14, -4, 39, 5, -40, 10, 10, -63, -55, 55, 21, -29, 30, -65, 46, 65, -82, 5, -15, 28, 10, 3, 58, -86, -48, 1, 82, 19, -104, 62, -4, -8, 58, -77, 20, 13, -63, 12, 42, -27, 48, 64, -36, -34, 18, 29, -81, -40, 12, -6, 79, 23, -90, 25, 49, -52, 28, 23, -35, 58, -51, -14, 51, -18, 43, -61, -1, 90, -53, -47, -29, 19, -3, 22, 96, -96, -32, 11, -45, 69, 4, -53, -17, 27, 61, 8, -2, -1, -58, -15, 31, 3, -30, -26, -12, 100, 24, -124, 79, 79, -61, -58, -10, 43, 75, -47, -28, 42, -60, 61, -24, -29, 6, -42, 0, 43, 78, -4, -45, -71, -20, 77, 21, -71, 52, 27, -60, -38, 39, -2, 21, 91, -65, -79, 44, 7, -13, -3, 27, 60, -78, 29, 27, -72, -13, 25, -5, -49, 24, 39, -29, 6, 5, -7, 47, 35, 24, -17, 19, -49, 0, 60, -72, -63, 71, 61, -55, -32, -32, -2, 1, 1, 5, 10, 42, -31, 42, 35, -61, -22, -38, 20, 73, -56, 36, 27, -112, 80, 8, -93, 31, -9, 59, 46, -73, 44, -4, 5, -12, -37, 3, -30, 79, -15, 3, 8, -27, 63, -71, -62, 18, -19, 48, 70, -49, -5, -15, -27, 52, -27, -7, 58, -14, -35, -8, 45, -14, -11, 52, -28, -47, 35, 51, 27, -71, -32, 35, 13, 8, -58, 64, 4, -53, 24, -41, 30, -3, -57, 4, 25, 27, -2, -24, 12, 70, -34, -51, 78, -51, 0, 48, -98, 56, -10, -66, 74, 43, -31, -20, 52, 41, -69, -29, -11, 43, 20, 0, 43, -39, 23, -22, -99, 20, 37, 25, -41, 27, -2, -99, 92, 86, -72, 17, 27, -60, -28, -31, 96, 26, -51, 58, -23, -100, 6, 57, 34, 25, -32, -14, 7, -8, -56, 0, 99, -17, -61, -32, 8, 21, -18, -7, -3, 43, -12, 3, 97, -66, -5, 81, -19, -37, 26, -44, -24, 10, 12, 30, -75, 5, -5, 24, 83, -61, -63, 69, 32, -38, 40, -69, 4, 19, -76, 2, 40, 22, 6, 27, -24, 20, -6, -21, -15, 0, 26, 49, 10, -49, -29, 48, 42, -37, -14, 10, 34, -81, -28, 68, -8, -9, 1, -1, -13, 38, 0, -62, -29, 4, 54, 36, 25, -43, -73, 10, 42, 62, -51, -30, 9, 26, 17, -59, 12, 1, -46, 26, 11, 37, -18, -85, 25, 71, 4, 12, 20, -88, -48, 80, 6, 5, 27, -56, -38, 41, 41, 9, -6, 12, -24, 2, 39, -7, -32, -60, -5, 10, 56, 7, -61, 37, 32, -38, 18, -54, -1, 15, -47, 40, 74, -20, -42, -7, 30, 27, -77, -11, 32, 26, -21, 11, 29, 15, 2, -1, -41, -3, 7, 12, 5, -54, 49, 36, -65, -63, 95, 21, -68, 68, -30, -80, 47, 11, 25, -53, 43, 57, -70, -9, -28, 44, -24, 3, 60, -21, 3, 18, -26, 11, 31, -23, -19, -29, 15, 2, 18, 0, -65, -27, 44, -4, -18, 74, 10, 4, 41, -39, -26, -27, 37, 58, -119, 36, 59, -59, 36, -49, -19, 5, -35, -6, 74, 34, -34, -20, 58, -20, -20, -6, -49, 26, -31, 47, 74, 1, -39, 22, -18, -69, -1, -2, 78, -7, -74, 28, 43, 47, -22, -61, -56, 53, 18, 22, -24, 2, 20, -76, -15, 89, 7, -62, 3, -5, 4, -32, -3, 56, 82, -44, 10, -34, -22, 87, -44, -75, 3, 3, 60, 71, -80, 30, 10, -40, 49, -15, -12, -63, 19, 82, -108, 51, 18, -105, 47, 1, -23, 21, 82, -57, 0, 92, -95, 0, 43, -23, 12, 22, 2, -15, 2, -58, 13, -7, 15, 41, -21, 2, -23, 20, -49, 6, 49, -53, 15, 76, -51, 9, 6, -82, 86, 2, -100, -5, 92, 31, -28, 15, -37, -6, 0, -52, 24, 105, -60, -45, 34, 25, 65, -99, -40, 13, -3, 98, -37, -76, 60, 43, -65, -65, 97, -3, -83, 108, -11, -77, 28, 70, 25, -6, -24, -89, 72, 0, -94, 12, 41, 54, -71, -2, 64, -24, 11, -24, -37, 82, 7, -86, 17, 51, -41, -17, 48, 8, -43, 39, 40, -14, 19, -26, 1, -28, -3, 53, -47, 15, 63, -95, -41, 100, 8, -87, -9, 22, -23, 64, -27, 8, -24, -10, 59, -66, -3, -24, 54, 62, -98, 5, 44, 31, -21, -65, 26, -24, -36, 89, -4, -104, 105, 61, -111, 5, 87, -34, 27, -27, -60, 21, -41, 8, 102, -3, -34, -17, -6, 18, 22, 30, -90, -19, 60, -21, 6, 66, -45, -5, 43, -53, 23, 36, -102, 46, 15, -14, 35, -66, -40, 63, 44, -82, -17, 36, 26, 35, 19, -69, -35, 40, 49, -34, 23, -1, -36, 51, -46, -56, 21, 87, 2, -64, 11, 35, -43, 30, 20, -9, -34, -20, 56, -12, 8, 38, -66, -55, 74, 39, -12, -73, -6, 35, 3, -5, 35, -10, -68, -8, 19, 66, -32, -64, 1, 66, 60, -42, 8, -11, -32, -27, -29, 3, 48, 92, -93, 5, 35, -18, 44, 20, -69, -74, 57, 21, 36, -39, 11, 77, -49, -54, 30, 26, -30, 32, 4, -63, 11, -8, 18, 70, -60, 10, -18, -102, 103, -22, 20, 4, -20, 88, -111, 45, -10, -51, 70, 0, 43, -32, -8, -9, 22, 22, -94, 14, 31, 0, 63, -68, -98, 103, -21, -43, 94, -60, -9, 60, -57, 5, 60, -53, -40, 87, -32, -48, 35, 32, -24, -34, 2, 54, 66, -86, -10, -29, 40, -1, -25, 107, -93, 9, 73, -90, -12, 28, -14, -43, 70, 37, -35, 19, 3, -55, -28, 87, -15, 7, 9, -20, -28, 11, 55, -76, -51, 22, -12, 79, -1, -14, 73, -74, 17, 7, -28, -14, 17, 68, -62, 0, -7, 34, -5, -1, -18, -32, 85, -38, -2, -17, -59, 80, -25, -23, 119, -102, 22, -7, 1, 18, -24, 73, -57, 17, -28, -86, 89, 78, -15, -62, -11, -1, -54, 97, -26, -70, 68, 35, 23, -48, -71, -12, 7, -7, 77, -7, -85, 96, -15, -79, 94, 71, -6, -53, -2, -39, -25, 65, 41, -43, 0, 28, -46, -25, -6, 38, 11, -51, -13, 36, -10, 6, 3, -3, 22, -31, -10, 48, 43, -27, -10, 46, -47, 0, -7, -69, 54, 53, -5, 7, -80, 15, 15, -35, 77, 8, -82, -21, 68, -7, -4, 58, 18, -94, -34, 40, -36, 44, 90, -82, -72, 80, 51, -9, -27, -69, 53, 3, -11, 48, -14, 42, -46, -89, 28, 7, 11, 34, -9, -29, 46, 3, -83, 69, -4, -4, -23, -18, 61, -68, 14, 75, 10, -24, -21, -18, 15, 8, -14, 25, -54, -3, 45, -11, 21, -60, 20, 30, -23, 8, 0, 22, 8, -60, -19, 8, 23, 45, -7, -24, -2, 25, -63, 32, -22, 29, -7, -5, 39, -20, 20, -19, -2, -46, -5, -7, 5, -5, 4, 95, 0, -85, 26, 9, -31, -14, 18, -8, 30, 10, -32, 28, 12, 40, -75, 13, 66, -82, 30, -8, -80, 29, 64, 8, -38, 60, 0, -10, -37, -86, 82, 51, -55, -20, 61, 22, -35, -31, 36, -8, -19, 2, 18, 17, -71, -30, 7, 85, 0, -93, 78, 28, -62, 34, 55, -81, -15, 57, -3, 34, -26, -6, -28, 48, -28, -76, 72, 22, 3, -3, -74, -14, 88, 32, 4, -95, 24, 9, -10, 23, -82, 71, 27, -10, -7, -27, 38, -26, -79, 37, 96, 4, -82, -19, 54, -24, 19, -8, 22, 22, -32, 60, 2, -35, 5, 4, -18, 6, 17, -29, 29, -43, -71, 60, 30, 34, -76, -39, 115, -45, -111, 103, 69, -83, -26, 10, 26, -32, 5, 47, -14, -4, -4, 10, -42, 2, -6, 51, 10, -102, 44, 18, -53, 65, 57, 2, -14, 0, -14, -10, -46, -12, 70, 0, 36, -71, -74, 61, -15, 23, 87, -7, -72, -7, 3, -24, 81, -4, -60, -17, 5, 73, -22, -23, 47, -59, 0, 31, -60, -13, 0, -13, 62, 48, 9, -14, -2, -41, -87, 94, 92, -112, -2, 17, -27, 90, -6, -34, -4, -68, 37, 91, 7, -76, -23, 54, -24, -23, -46, 29, 52, -68, 40, 0, 3, 47, -13, 2, -19, 35, -14, -40, 56, -41, -21, 51, -65, -2, -6, 21, 19, 28, 23, -64, -25, 0, -29, 41, 63, -78, -13, 5, -34, 111, 4, -117, 49, 99, -5, -79, 44, -23, -7, 79, -63, -5, -4, -14, 77, -9, -83, 7, 18, 28, 32, -5, -83, 24, 35, -40, 61, -5, -13, -60, -3, 99, -70, -63, 89, 32, -31, 0, 32, -20, -32, -6, -49, 52, 90, -85, -46, 6, 12, 60, 36, -41, -59, 87, -41, -23, 64, -92, -2, 25, -43, -3, -5, 1, 22, 62, 35, 9, -29, -21, -10, 27, 61, -62, -6, 38, -11, -80, 46, 3, -18, 81, -41, -53, 32, 52, -76, -34, 74, 9, -29, 35, 4, -17, -56, -61, 43, 87, -51, -95, 65, 46, -64, -2, 96, 35, -75, -25, 90, -53, -23, 93, -85, -41, 37, -49, -8, 49, 26, -46, -27, 20, -35, 68, 96, -114, 30, 26, -4, -23, -69, 63, 0, -21, 58, 7, -79, 3, -17, -9, 39, 72, -48, -18, 29, -35, 42, 18, -72, -41, 82, -10, -41, 68, -32, -58, 88, -26, -31, 88, -73, 36, 12, -52, 35, -38, -42, 44, 57, -85, 61, -15, 9, 9, -35, 41, -24, 8, 35, 14, -29, 5, 22, -48, -59, 103, 0, -82, -9, -31, 92, 25, -104, -1, 85, 18, -63, 68, -47, -5, 96, -9, 0, 14, -93, -13, 30, -5, -4, -43, 11, 52, 73, -75, -89, 35, 5, 3, 44, -27, -2, 22, -1, 3, 18, -6, -70, -22, 34, -4, -29, 21, -13, 79, 15, -104, 65, 23, 6, 37, 2, -74, 0, 75, -61, 26, -23, -31, 28, 0, 51, 25, -65, -41, 28, 41, 39, -40, -69, -36, 68, -9, -36, 77, -42, -21, 85, 22, -87, -2, 78, -87, -73, 59, 77, -21, -48, 80, -56, -19, 80, -6, 26, -102, -26, 54, -57, -5, 106, -37, -40, 61, -27, -53, 4, 40, 36, -20, -49, 80, -22, -100, 108, -10, -38, 76, -11, -68, 21, 66, -90, -8, 60, 24, 2, -75, -29, 54, 30, -58, 39, -10, 3, 9, -64, 7, 52, -28, -11, 4, 28, 76, -97, 28, 64, -4, -8, -36, -54, 10, 8, -29, -20, 72, -2, -19, -3, -30, 36, 1, 46, -60, 14, 48, -48, -48, 56, 1, -78, 44, 4, -24, -15, 44, -20, 48, 39, -29, 12, -12, -15, -1, 69, -38, -17, -24, -59, 68, 34, -23, -14, -31, 48, -24, 17, -1, -73, 77, -20, -39, 97, -11, -62, 81, 27, -62, 40, -24, -70, 31, 48, 25, -79, 30, -13, -8, 97, -73, -27, 17, 14, 44, -15, -25, -69, 2, 61, -29, -52, 43, 43, 20, 53, -111, 10, 80, -60, 29, 30, 3, -49, -5, 25, -18, 4, 10, -6, -12, -40, -36, 6, -22, -12, 82, 40, -82, 0, -8, 0, 35, 11, 65, -38, -26, -22, -26, 28, 27, 4, -47, 31, 63, -54, -52, 44, 60, -40, -71, 48, 8, -13, 34, -15, -3, 5, 25, 25, -20, 38, -64, -78, 71, -23, -2, 23, -64, 87, 26, -11, -22, -2, 39, -70, -53, 74, 86, -106, -52, 14, 30, 44, 1, -22, -59, -1, 68, 76, -88, -37, 115, -66, -1, 51, -65, -2, 48, 3, -30, -10, -11, 57, -10, -85, -13, 44, -6, -58, 54, 26, -41, -22, 72, 70, -71, 35, -25, -90, 113, -26, -13, 94, -70, 5, 8, 0, 0, -54, 26, -54, 51, -9, 4, 39, -93, -5, 62, 10, -63, 6, 36, 2, -18, 21, -40, 45, 30, -64, -20, 7, 42, -35, -28, 87, 57, -21, -2, -32, -52, 0, 25, -25, -5, 35, -9, 11, 29, -58, 22, 75, -53, -27, -32, 41, 79, -74, 0, 0, -27, 68, 9, -94, 31, 89, -8, 0, -24, 8, -37, -76, -10, 81, -12, -15, 4, 0, -4, 10, 76, -96, 0, 22, -37, 77, -46, -43, 3, 42, 44, -25, 22, -58, 12, 52, -82, 27, 26, 6, 17, -28, 43, 3, -37, -60, -12, 58, 28, -18, -18, -8, 20, -41, -5, 98, 12, -28, -61, 38, 11, -17, 37, -103, 58, 27, -49, -21, 34, 89, -14, -38, -32, 46, -35, -91, 79, 41, -29, -4, 45, -49, -15, 66, -91, 2, 27, 57, -49, -28, 95, -42, -23, 0, -6, 8, 27, -56, -12, 62, 29, -5, -91, 21, 18, -37, 46, -37, 29, 12, -42, 75, -38, -31, 6, -17, 58, 39, -71, 27, 27, -87, -10, 93, 2, -18, 13, -83, 59, -22, -17, 90, -54, 30, -24, -10, -5, -4, 86, -90, -77, 44, 75, -26, 11, -27, -19, 68, 6, -68, -13, 36, -66, 88, -4, -39, 68, -15, 13, -8, -15, 15, -31, -44, 23, 35, 32, 18, -54, 5, 37, -21, -59, 0, 87, -71, -26, 66, -1, -17, -2, -12, -6, 65, -61, 10, 45, -107, 20, 37, -4, 6, -78, 76, 47, -54, 24, -9, -17, -32, -2, 0, 37, 28, 4, 10, -22, -2, -34, -20, 68, 53, -31, -25, 4, 35, -15, -59, -46, -17, 68, 40, -32, 13, 3, 32, -19, -82, 25, 52, -23, 1, 76, -78, -59, 77, 42, -81, -35, 7, 8, 32, -52, 0, -15, 69, 12, -29, 11, -56, 64, 55, 6, -59, -22, 32, -46, 49, 39, -21, 11, -77, 3, 62, -45, -55, 30, -1, -45, 88, -17, -11, 11, -68, 95, -8, -85, -3, 72, 13, -59, 48, -19, -52, 77, 46, -18, -60, 5, 19, 30, -4, -57, 37, 36, 10, -18, -42, 9, 68, -91, 18, 53, -82, -25, 11, 24, -21, 10, -12, -8, 64, 12, -29, 32, -1, -72, 15, 27, 21, 35, -29, -72, -21, 95, 54, -10, -11, -81, 19, 32, -57, 15, 64, -26, -7, -32, -2, 82, -46, 6, -17, -72, 19, 43, 52, -3, -6, -23, -66, 36, -10, -4, 54, -31, 1, 14, -20, -34, 48, -21, -22, 105, -5, -48, -11, -12, 26, -15, -40, -15, 78, 29, -87, 9, -14, -35, 94, 65, -58, -59, -7, 41, 25, 22, 30, -62, -51, 10, -7, 86, -9, -117, 78, 95, -56, -47, -4, -26, 23, 42, -40, -6, 74, -14, -20, 58, -30, -17, 36, -91, 34, 3, -45, 59, 25, -13, -4, -25, -4, 9, -49, -12, 3, 8, 61, 59, -42, -32, -56, -18, 100, -8, -21, 63, -6, -22, 7, -13, -39, 20, 8, -28, 27, -37, 30, 55, -53, 27, 28, -36, -76, -19, 40, 18, -10, 11, -11, -53, 70, 19, -70, 58, 31, -72, 9, 25, 15, -2, 9, -1, -94, 20, 61, 21, -18, 3, -13, -51, 28, -5, 6, 43, -23, -63, 63, 75, -53, -61, 44, 13, -42, -2, -40, -7, 13, 58, 17, -59, -34, 27, 29, -37, 26, 92, 4, -81, 5, -12, -19, 13, -17, -12, 36, 73, -80, 11, 37, -23, 61, -30, -97, 20, 55, -46, -7, 73, 10, 9, 11, -3, -49, -70, 68, 86, -91, -11, 4, 3, 65, -38, 41, -63, -27, 78, -14, 24, -24, -68, 23, 13, -7, 17, 36, -64, -6, 25, 5, 26, -77, 40, 1, -39, 83, -40, -40, -8, 34, 54, -3, 10, -74, 37, 55, -102, 5, 40, 34, -42, -25, 59, -30, -11, -36, 8, 12, 46, 35, -70, -37, 69, 58, -32, -57, 27, 36, -8, 20, -19, -47, 39, -34, -9, 78, -112, 24, 58, -69, 60, 14, -74, 7, -11, 0, 63, -3, -76, 21, 27, -36, -13, -11, 23, 37, 43, -60, -15, 55, -42, -35, 9, -26, 44, -17, 30, 65, -109, 3, -5, 63, -3, -78, 74, -20, -52, 2, 87, -18, -86, 7, 57, -10, -23, 80, 46, -71, -70, 31, 73, -22, -2, -29, -26, 40, -47, 7, 86, -42, -14, 104, -91, 2, 22, -18, -17, -27, -12, 47, 63, -99, -31, 8, 3, 29, 90, -61, -17, 18, -29, 54, -5, -30, 24, -29, -12, 87, -25, -15, -45, -19, 61, -21, -35, 63, 72, -56, -54, -29, -8, 99, -37, -61, 109, -36, -6, 85, -77, -3, -34, 29, 25, -41, 24, -85, 64, -11, 4, 41, -52, 71, 20, -79, -41, 3, -15, 8, 39, 21, -43, 56, 5, -59, 15, -20, 38, 6, -47, -14, -22, 32, -3, -15, 106, -4, -75, 55, 2, -46, -39, 85, 1, -15, 7, -62, 100, -32, -28, 28, -13, 62, -51, 17, 0, -35, -1, 17, 86, -73, 4, 62, -20, -91, -43, 85, -7, -3, 7, -5, 58, -32, -8, -29, -51, 86, 18, -61, -34, -10, 57, 63, -61, -82, 81, 27, -6, -31, -43, 78, 5, -41, 29, -11, -23, -11, -60, 81, 72, -51, -9, 14, 48, -43, -13, 21, -70, 7, 48, -14, -1, 15, -63, 51, 20, 17, -11, -74, -14, 30, 93, -8, -95, 11, 89, -29, -21, 51, -39, -37, -2, 57, -21, -62, 15, 54, 46, -53, -24, -18, 64, -52, 1, 2, -3, 22, 20, -15, -51, 4, 15, 44, -28, 53, -58, -25, 19, 32, 2, -18, -3, -1, 39, -25, -62, 56, 27, -17, 2, 0, -9, -64, 60, 78, -62, -29, 10, -44, 43, 51, -38, -28, -20, 65, 0, -75, 38, 21, -41, 39, 3, -44, 41, 19, 39, -22, -12, -24, -19, -10, -45, 61, 13, 19, 27, -27, -10, 13, 61, -81, -23, 22, -21, 72, -46, 2, -4, -8, 22, -44, 34, -1, 42, -37, -68, 80, 47, -81, -54, 30, -2, -5, 70, 32, -79, 7, 3, 19, 23, -45, -38, -21, 66, 49, -62, -66, 54, 22, 14, 55, 0, -41, -35, 38, 31, -102, 9, 78, -72, -62, 90, 37, -73, 73, -42, -15, 55, -39, 25, -32, -82, 76, 34, -13, 19, -30, 49, -40, -97, 89, -11, 15, 25, -45, 80, -80, -10, 69, -21, 28, 3, -21, -25, -44, 24, 41, -61, -26, 6, 52, 27, -73, 20, 61, 43, -75, -57, 95, -27, -39, 48, -17, -3, -38, -38, 54, -30, 63, -10, -27, 91, -8, -26, -48, -30, -23, 86, -2, -48, -18, 51, 89, -94, -18, 58, -51, 15, 3, -89, 103, 52, -39, -2, -64, 32, 49, -34, 26, 0, -24, 20, -23, -8, -29, 19, 51, -52, -4, 47, 8, -25, 11, -14, 11, -7, -88, 76, 95, -82, -99, 85, 77, -28, -29, -74, 5, 106, 3, -77, 18, -23, 53, -25, -28, 22, -7, 20, -30, 7, -41, -18, 72, 58, -31, -22, 48, 10, -59, 34, 37, -48, 7, 24, -55, -44, 39, 60, -49, -43, -17, 55, 46, -96, 53, 14, -75, 46, 14, 8, 31, -27, 9, 12, -60, -2, -12, -9, -12, 42, 0, 23, 13, -102, 51, 44, -35, -18, -2, 25, 25, -17, -28, 71, 15, -86, -22, 53, 46, -7, -26, -12, -13, -14, -19, 14, 74, -52, 6, 61, -13, 30, -27, 18, -53, -89, 68, 1, -14, 44, 24, 31, -64, -92, 104, 38, -69, -30, 6, -22, 49, 70, -35, -52, -59, 58, 53, -7, 28, -31, -39, 34, -2, -63, 35, 30, -38, -28, 35, 56, 12, -25, -25, 60, -7, -31, -11, 34, 24, -5, -76, -13, 64, -20, 21, 4, -52, -17, 19, -46, 42, 69, -7, -72, 26, 22, -40, -11, -4, -3, 42, 7, -31, 40, -46, -15, -15, 56, -1, 9, 51, -81, 20, -21, 34, 15, -13, -14, 0, 3, -61, 44, 51, 40, -29, -11, -24, -69, 65, 57, -71, 0, 63, 28, -75, -69, 13, -2, 76, 11, -79, 13, 43, 25, -6, -9, -46, -21, 63, 42, -18, -88, -2, 28, 62, -32, -90, 40, -12, 64, 76, -60, -28, 52, -34, 8, -38, -18, 4, 37, -4, -75, 53, 35, -25, -66, 27, 14, 22, -17, -30, 2, -15, 56, 35, -63, 25, 57, -48, 32, 30, -63, -7, 2, -32, 73, -11, -70, 55, -6, -31, 28, 30, 19, -44, 5, 62, -18, -66, -26, 75, -9, -23, -30, -41, 11, -5, 75, 47, -31, 15, -14, -71, -12, 76, 8, -73, 66, 48, -20, -27, -75, 28, -18, 38, 74, -13, 11, -36, -61, -13, 18, 21, 54, -32, -18, 64, -17, -36, 19, -27, -20, -14, -7, 56, 41, 0, 4, 18, -42, 5, -36, -3, 13, -55, 57, -25, -44, 47, 28, -15, 32, -42, -85, 88, 10, 7, 41, -94, -6, 38, -30, 66, 1, -19, 31, -48, 0, 35, -29, -40, 17, 47, -64, 34, -7, -6, 7, -51, 43, 9, 66, -58, -5, -20, 29, 5, -11, 71, -91, 6, -27, 11, 46, -25, 19, -57, 60, -3, -19, 29, -45, 23, -59, 26, 32, -66, 22, 19, -4, 42, 52, -28, -106, 45, 40, 11, 49, -61, -7, -17, -75, 55, 82, -27, -58, -10, 49, -22, -12, 28, 7, -54, 29, 59, -27, -47, 13, -7, -28, 9, 35, 24, -42, 62, -44, -89, 77, 93, -39, -39, -37, 17, -7, 48, -11, -64, 40, 14, 25, 23, -42, -78, 79, 75, -18, -39, -62, -1, 43, -4, 10, -31, 41, -8, -104, 111, -11, -25, 92, -27, -65, 55, -11, -75, 108, -47, -4, 11, -8, 42, -99, 62, 51, -18, 47, -60, -34, -36, 27, 98, -38, -49, -24, 0, 27, -13, -21, 39, -19, -41, 9, 26, -6, -23, 88, -35, -44, 80, -26, -29, -13, 10, 8, 37, 12, -55, -20, 65, 20, -103, 56, 90, -44, -78, 5, -15, -3, 75, 1, -18, 30, 30, -83, -63, 6, 94, -8, -37, 62, -12, -70, 49, -3, -62, 89, -12, 15, -46, -34, 35, -39, 24, -4, 29, 35, -22, 34, -58, -36, 32, 30, -3, -66, 59, 19, -56, 43, 29, -75, -5, 17, -30, 22, -9, 44, -24, 1, 60, -73, -29, 73, -1, -5, -22, -61, 28, 44, 62, -30, -81, 7, 0, 4, 32, 40, 24, -3, -7, -36, -54, -36, 71, 5, -32, 63, 47, -38, -24, -4, -1, 56, -42, -89, 48, 22, -58, 55, 91, -87, -64, 7, 9, 26, -7, 66, -23, -73, 60, 58, -17, -15, 42, -39, -103, 32, 3, 37, 82, -19, -56, -7, 35, -12, 18, -47, 9, 93, -108, 12, 6, -83, 115, -4, -32, 15, -51, 53, 53, -104, 23, 32, -6, 47, -29, 26, -56, -2, 85, -89, -1, 27, -95, 35, -6, 17, 77, 3, -2, -6, 15, 1, -68, 14, 18, -99, 10, 55, 68, -71, -21, 89, -41, -5, 22, -44, -3, 77, -48, -29, 11, -48, -22, 7, 74, -30, -63, 63, -28, 45, 34, -10, 46, -35, 28, -71, 1, 14, -12, 69, -58, -10, 21, 35, -17, -69, 10, -21, -11, 55, 41, -19, 8, 13, 10, -29, 5, -54, 10, 90, -9, -43, -12, 55, -77, -7, 97, -75, -103, 86, 81, -49, -36, 15, -13, 36, 38, -24, 36, -64, -58, 73, 24, -48, -20, 35, 32, -37, -18, 68, -62, -6, 20, -74, 29, 35, 30, -6, -40, 60, -34, -45, 9, 20, 59, -5, -31, 5, -7, -19, 29, 46, -58, -30, -5, 28, 4, -81, -5, 75, 75, -68, -19, -15, -30, 98, 18, -88, 0, 0, -51, 58, 42, -41, -5, -10, 64, 48, -4, -31, -62, 48, -9, -8, -5, -11, 24, -23, 15, 15, -36, -19, 61, 31, -35, -58, 40, -19, -35, 19, -37, 28, 57, 5, 8, -64, 17, 73, -20, 32, -71, -59, 59, 10, 21, 53, -92, -43, 29, 14, 62, -6, -94, 32, 24, -38, 65, 40, -32, -56, -52, 40, 58, 6, -41, -47, 73, -27, -81, 57, 94, -64, 0, 41, -34, 46, -42, 9, -23, -11, 49, -73, -18, 43, 49, 6, -82, 27, 45, -4, -53, -2, 37, 3, 3, -7, -18, -56, 78, -11, 3, 61, -58, 23, -9, -68, 43, 61, -80, 21, 48, -30, -49, 27, 35, -112, 37, 41, 25, -27, -71, 85, 57, -35, -1, -27, -41, 68, 27, -74, -35, 53, -38, 20, 55, -47, -23, -13, 12, 7, -12, 62, -22, -62, 94, -9, -38, -5, 54, -15, -32, 6, -44, 22, 83, -68, -3, 63, -112, 24, 78, -30, -56, 65, -13, -1, 15, -36, -11, 6, 82, -28, -17, -30, -70, 54, 46, 3, -60, -7, 98, -6, -2, -34, -72, 78, 6, -75, 11, 6, 61, -45, 0, 3, 19, -11, 2, 35, -49, -9, 42, 34, -37, 25, -22, 26, -34, -62, 29, -7, 43, -5, 8, 40, -43, -39, -14, 78, -26, -4, 0, -77, 61, 89, -72, -31, 97, -72, 3, 48, -81, 43, 80, -96, -41, 61, 19, 12, 1, -61, 25, 44, -70, 57, -30, -88, -3, 44, 79, -27, -66, 77, 25, -119, 55, 63, -37, 15, 14, -13, -47, -42, 28, 12, -46, 77, 74, -119, 0, 75, -71, 27, -14, -4, 62, -64, 20, 34, 5, -13, 25, -43, -48, 52, -52, 7, -17, 46, 0, 1, 35, -70, 71, 39, -32, -68, 24, 38, -76, 26, -20, -9, 29, -34, -12, 71, 10, 5, 14, -75, 14, 18, -5, -54, 49, 57, -72, 56, -7, -47, 55, 1, 15, 12, -44, -19, 52, -19, -90, -21, 97, -20, -30, 17, -53, 70, 62, -20, -13, -36, 39, -24, -17, 35, -78, 34, 68, -14, -23, -28, -41, 5, 86, -23, -92, 41, 47, 54, 0, -19, -57, -15, 72, 0, 1, -70, -21, 59, 22, -56, 26, 60, -81, 12, 69, -26, -65, 53, -42, -1, 113, -83, -82, 87, 3, -62, -7, 77, -11, -7, 58, -73, -2, 15, -45, -24, 37, 24, 37, -53, -11, 66, -14, 39, -36, -31, 11, 8, -3, -28, 32, -25, -2, 61, -69, 4, 107, -80, -6, 3, -66, 28, 24, 22, 24, -20, 18, -29, -88, 57, 4, 13, -10, 11, 52, -44, -20, 62, -35, -23, 32, -4, -47, 31, 56, -120, 61, 27, -62, 31, 11, -14, 34, 59, -82, -29, 37, 23, 28, -46, -29, 56, -35, -39, 70, 13, -63, -63, 80, -10, 26, -19, -15, 112, -99, -69, 104, 48, -39, -49, -9, -30, 45, 28, -103, 75, 83, -65, 14, -1, 17, -17, -53, -15, 54, -5, -21, 105, -72, -32, 2, -45, 58, -11, -66, 70, 28, -73, 11, 100, -36, 3, -20, -80, 28, -11, -23, 94, 36, -13, 3, -34, -30, 35, 60, -89, -58, 60, -8, -17, 7, -26, 51, 46, -40, 5, 5, -11, 43, 14, -1, -82, 18, 68, -71, 26, 57, -75, 27, 0, -66, 7, 55, 13, -66, 6, 39, -36, 46, 30, -54, 53, 23, -93, 10, -14, 0, 106, -25, -47, 29, -28, -15, 28, 15, 45, -60, -15, -5, -54, 74, 17, -43, 20, 29, 20, -85, -41, 97, 48, -8, -44, 11, 13, -27, 0, -1, -3, -8, -7, -49, 2, 54, 21, 29, -19, -22, -7, -59, 60, 49, -96, -8, 4, 35, 0, 5, 61, -43, 14, 15, -31, -30, 28, -19, -57, 8, 69, 28, 2, -51, 0, 1, 2, 43, -82, 7, -1, 0, 60, -52, -58, 76, 26, -52, -1, 46, -25, -53, 5, 80, 54, -27, -38, -28, 63, -7, -19, 42, -68, -14, 80, 20, -13, -4, -26, -74, -21, 62, 18, 20, 10, -20, 5, -75, 40, 91, -27, -70, -77, 110, -14, -21, 82, -54, -27, 30, -40, -46, 54, -19, 48, 23, -88, 57, -3, -24, 72, -23, -49, 0, -6, 74, -42, -2, 21, -113, 91, 82, -94, 13, 83, -89, 14, 28, -9, -10, -72, 64, 29, -15, -45, -11, 5, -22, 22, 2, -21, -40, 92, 14, -40, 0, -25, 51, -25, -26, 72, -46, -53, 85, 78, -80, -91, 93, 34, 13, -51, -9, 74, -23, -26, 29, -34, -21, 7, -12, -17, -35, 60, 49, 3, -70, -41, -20, 70, 21, -44, 31, -26, 34, 6, -59, 62, 24, -77, 9, 36, -19, 0, 0, -22, -27, 11, 35, 39, 22, -88, 23, 97, -29, -13, -10, 11, 32, -34, -7, -36, -56, 0, 27, 70, -14, -4, 20, 6, 48, -83, -43, 27, 5, 49, -14, 0, -30, -70, 40, 78, -46, -45, 62, 56, -60, -60, 89, -31, -89, 60, 23, -53, 37, 73, -74, -68, 66, 57, -60, -17, 85, 6, -99, 4, 52, -4, -14, 1, 37, 24, -32, 10, -1, -81, 70, 24, -28, 26, -5, 12, -27, -71, -17, -11, 94, -3, -76, 52, 48, -2, -78, 47, 0, -68, 31, 32, 40, 14, -55, -12, 39, 20, -2, -72, -36, 41, 62, -64, -38, 60, 38, 21, -10, -69, -79, 83, 13, -44, 26, -44, 62, 35, 5, -48, -9, 35, -18, 52, -61, -49, 13, 88, -29, -96, 18, 22, 38, 59, -20, -93, 29, 13, 41, -2, -55, -11, -52, 73, 30, -46, 53, -19, 10, 56, -72, 22, -20, -68, 51, 9, -27, 69, -10, -57, 86, -18, -13, 31, -48, -34, 29, 72, -19, -18, -19, -75, 58, 19, 0, -22, -5, 49, -44, 29, -30, 19, 29, -51, -44, 58, 71, -71, 17, 55, 2, -10, -53, 10, -4, 10, -21, -85, 85, 44, 11, -68, -6, 68, -49, -6, 42, -34, -69, 0, 83, 10, -90, 2, 71, -23, -47, 28, 35, -32, -23, 40, 41, 35, -59, -48, 45, 5, -20, 18, -37, -11, 59, -43, -53, 11, 39, 81, -44, -6, -9, -49, 4, -8, 42, 56, -31, 15, -25, 1, 91, -52, -46, 44, -20, 3, -2, -86, 10, 66, 21, -25, -30, -29, 41, 2, -19, -5, -26, 48, 77, -57, 0, 79, -44, -46, 20, 55, -54, -5, 80, -76, -36, 34, -53, 56, 17, -75, 82, 24, -97, 17, -1, -39, 77, 17, -10, -52, 10, 72, -7, -2, -76, 14, 51, -9, -29, -36, 44, 24, -40, -5, 59, 31, -83, -78, 88, 19, -39, 39, 45, -5, -58, -45, -22, -3, 61, 55, -55, -14, 34, -39, -38, 49, 65, 11, -49, -54, -25, 85, 59, -65, -9, 31, -34, -6, 64, -58, -74, 23, 88, -28, -91, 31, 13, -21, 9, 78, 30, -25, -26, -45, 46, 20, 3, 23, -57, -46, 56, 29, -71, 6, 72, 28, -71, -53, 42, -27, -19, 56, -1, -40, 26, 19, -29, 44, -4, 0, 30, -64, -24, 90, 0, -89, 25, 4, 22, 57, -42, -8, -26, 18, -2, -64, 47, 14, -24, 70, -11, -22, 14, -17, 69, -70, -83, 38, 60, 21, -70, -18, 65, 14, -37, -42, 37, 75, -38, -29, 40, -58, -59, 105, 47, -60, -45, -17, 63, 38, -60, -34, 13, 64, -47, -49, 108, -45, -7, 56, -4, -58, -73, 63, 44, -20, 21, -7, -38, 3, -38, -15, 34, 13, -20, -26, 66, 19, -44, 43, -54, 8, 96, -39, -36, 45, 43, -41, -89, 55, -8, 0, 86, -82, -21, 14, 30, -25, 9, -4, -43, 88, -45, 13, -8, -66, 98, 31, -24, -34, -39, 54, -28, -53, 13, 44, -4, -53, 3, -3, 94, -4, -91, 66, 21, -3, -28, -35, -6, -41, 52, 40, 23, 31, -60, 34, -12, -73, 69, 46, 2, -78, -7, 86, -43, 9, 17, -25, -43, 18, -7, -63, 14, -8, 94, 38, -102, -45, 114, -22, -85, 54, 39, -39, -28, 3, -27, 48, 19, 41, 6, -70, -17, 0, -4, 52, -11, 13, 24, -56, 34, -3, -4, 23, 7, 0, -51, 14, 66, -71, 19, -20, -14, 58, -61, -41, 38, 25, -15, 79, -25, -97, 9, 45, -9, 6, -11, 1, 20, -9, 57, 49, -105, -36, 73, 14, -58, 26, 29, 3, -19, -61, -14, 52, 83, -74, -74, 10, 59, 19, -41, 37, 31, -30, -28, 44, -26, -41, 44, -8, -28, -9, 42, -24, -43, -15, 102, 7, -103, 45, 12, -34, 71, -1, -66, 44, 31, -31, -53, -18, 97, 12, -93, 43, -20, -8, 64, -47, -24, -24, 55, 32, -29, -11, 7, 35, -27, 1, 39, 0, -64, -56, 78, 95, -59, -76, 28, 85, -22, -26, -20, -13, -15, 0, 4, -36, -4, 48, 27, -54, 48, -29, 0, 13, -39, 12, 27, 42, 10, -19, -70, 56, 32, -100, 42, 81, -66, -39, 56, 45, -92, 38, 32, -108, 40, 17, -29, 10, 69, -3, -21, 3, -10, -20, -4, 59, -8, -65, 10, 1, 1, 57, -74, 35, 66, -29, 6, 19, -51, -49, 66, -29, -30, 80, -27, 8, -12, -37, 39, -60, -17, -1, 34, 60, -20, -56, 7, 80, -37, 24, -28, -14, 80, -104, 42, 32, -111, 47, 28, -46, -21, 77, 34, -54, 45, 27, -24, -80, -7, 107, -49, -22, -7, 4, 38, -52, 60, 45, -61, -65, 68, 19, -78, 12, 53, -59, 24, 54, -9, -54, 3, 100, -91, -51, 66, -47, -19, 22, -38, 86, -6, -64, 61, -14, -56, 76, 66, -110, 35, 3, -66, 81, 0, -10, -14, -56, 63, -14, 0, 54, -72, 27, 18, -27, -44, 64, 37, -63, -24, 20, 21, -53, 70, 59, -46, -78, 46, 19, -78, 60, 1, -6, 7, 26, -21, -9, -3, -92, 87, 82, -36, -72, 0, 92, -11, -41, 44, 45, -86, -93, 69, 24, -35, 27, -24, 28, 59, -88, -62, 94, 60, -61, -2, -21, -34, 64, 60, -61, -3, 56, -69, -39, 71, 41, -60, -28, 19, -17, -2, 23, 5, -65, 48, 80, -39, -64, 19, 19, -65, 73, -20, 18, 7, -23, -1, -27, 65, -78, 46, 36, -20, -21, -3, 52, 15, -42, -88, 39, 30, 0, 41, 38, -46, -1, 28, -89, 46, 27, -71, 3, -36, 46, -1, -25, 23, -26, 60, 66, -83, 12, 10, -82, -6, -11, 61, 100, -78, -3, 25, -25, 15, -43, 10, 77, -43, -70, 12, -21, 48, 36, -40, 36, -29, -20, 10, -30, 86, -40, -52, 2, 64, 51, -100, 58, 36, -15, 43, -22, 1, -43, -23, -7, 22, -7, -60, 91, 8, -46, -20, -31, -12, 28, 96, -43, -78, -3, 36, 96, -66, 7, 6, -94, 56, 17, -37, -20, 25, -19, 73, 5, -61, 48, -1, -35, 15, 70, -59, -60, 23, 10, 0, -11, 63, -15, -55, 96, -43, 6, 77, -89, 14, 60, -51, -39, -31, 23, 30, -27, 29, -11, 0, -29, 14, 109, -69, -54, 69, -18, -3, -39, -7, 106, -54, -29, -22, 24, 39, -70, 58, -17, -22, 46, 44, -73, 7, 12, -48, 37, -14, -14, 4, 96, -48, -65, 95, -10, -8, 30, -5, -13, -11, 7, -22, -40, -45, 45, 77, -27, 0, 21, -24, -3, -42, 19, 36, -56, 35, -13, -20, 20, -31, 8, -17, 30, 52, -34, -70, 63, -7, -74, 29, 73, 26, -12, 32, 3, -61, 17, -2, -62, 18, 64, 24, -25, -5, -30, -60, 6, 46, 11, 6, 17, 19, 7, -42, -18, -29, 0, 25, -56, 39, 29, 38, -23, -74, 92, -46, -21, 88, -48, -59, -7, 15, 54, 57, 11, -88, 20, 14, -39, 31, 18, 2, -61, 28, 47, 9, 0, -38, -77, 76, -23, -45, 115, -49, -96, 74, 14, -7, 29, -30, 42, 0, 6, 4, -30, 18, 25, -10, -76, 5, 18, -55, -11, 47, 85, -74, -28, 85, -27, 5, 27, -27, -17, 8, 32, -5, -27, -42, 9, -20, 40, 27, 1, -40, -79, 81, 64, -52, -38, -9, 43, 69, -66, -56, 27, 14, -21, -1, -11, -26, 4, -3, 36, 76, 5, -21, -15, -23, 47, -29, -42, 90, -1, -41, 45, -59, -71, 111, -24, 1, -10, -65, 72, 7, -7, -32, 46, -34, -35, 36, -83, 86, 6, -25, 72, -78, -25, 29, 10, 0, 0, -7, -21, -1, 62, 1, -61, 15, -23, 51, -4, -32, -13, 44, 89, -24, -76, 22, 49, 1, -76, -7, 86, -72, -9, 23, -36, 54, 30, 0, -36, -59, -7, 28, 51, -76, 32, 99, -62, -77, 39, 42, -21, 25, -2, -23, -1, 30, -1, -60, 34, 30, -66, -11, 73, 11, 10, -52, -24, 62, -74, 28, 93, -83, -29, 31, -27, 0, 0, 22, 34, -73, -22, 11, 41, 65, -11, -49, 8, -17, 0, 22, -6, 44, 7, -20, -32, 15, 36, -56, -53, 97, -30, -68, 14, 26, 53, -12, -59, -35, 8, 62, -18, -31, 74, 43, -58, -29, 14, -70, 44, 104, -46, -51, 58, -18, -75, 26, -21, 54, 59, -72, 40, 25, -8, -57, -32, 43, 18, 0, -12, 51, -52, -10, 39, -89, 36, 68, -5, -81, 21, 57, -91, -21, 97, 56, -40, -65, -29, 72, -37, 29, 21, -111, 81, -10, -55, 27, 12, 75, 25, -90, 32, -6, -99, 53, -7, 48, -7, -13, 98, -97, -64, 116, -10, -78, 64, 57, -35, -74, 17, 60, -68, 20, 64, -10, 29, -82, -73, 65, -29, 39, 87, -104, -76, 96, 38, -81, 34, 49, -74, -1, 63, -27, -18, 52, 25, -68, 22, -11, -31, 21, 27, 34, -73, 3, 44, -65, 14, 61, -20, 7, 10, -46, 13, 44, -59, -57, 73, 65, -28, 20, -27, -55, -7, 63, -4, -94, 22, -3, -13, 80, 15, -73, 3, 52, 41, -86, 12, 55, -26, 12, -51, -13, 77, -37, -80, 19, 13, -7, -25, 8, -6, 38, 42, -12, -6, 39, 2, -7, 35, 7, -17, -39, -46, -15, 13, -25, 12, 3, 29, -10, -3, 93, -26, -37, 54, 2, -17, -39, -3, 69, -55, 11, -7, 9, -4, -12, 49, -4, 1, -29, 26, -19, -66, -38, 56, 39, -86, 70, 42, -36, -31, -49, 55, 27, 25, -1, -55, 6, 68, -59, -36, 14, 40, 66, -86, -49, 51, 72, -54, -59, 66, -49, 13, 90, -90, -14, 14, -41, 31, 39, 37, -25, 10, 1, -88, 57, -24, -27, 43, 23, 24, 3, -51, -23, 70, -28, -75, 10, 46, -42, 65, -18, -68, 79, 45, -23, -47, -47, 46, 72, -8, -4, -44, 24, -28, -19, 60, -53, -25, -10, -7, 0, -25, 32, 66, 24, 5, 11, -58, -40, -6, -13, 29, 36, -43, -9, 10, -5, 53, -52, -20, 44, 29, 44, -42, -87, 49, -4, -48, 116, -37, -31, 1, -41, -1, 68, -18, 5, 80, -77, -30, 52, 19, -2, -23, -1, -14, -11, -4, 15, 47, -27, -29, -10, 18, 15, 13, -64, 9, 100, -85, -4, 66, -82, -42, 44, 97, -64, -38, 66, -32, 39, 6, -98, 38, 70, -11, 27, -53, 6, 41, -5, -22, 12, -15, -5, 27, -3, -47, -73, 96, -23, -73, 32, 6, -29, 79, -7, -74, 42, 34, 26, -27, -71, 39, 97, 0, -61, 31, -30, -58, 75, -59, 34, 65, -75, 52, -19, -79, 92, 20, -90, -42, 57, 31, -57, 51, 0, -64, 88, 18, -5, 3, -12, 55, -71, -4, 53, -20, 6, 22, -57, -34, -14, -20, 8, 21, 11, -31, 80, -30, -10, 99, -74, -40, 17, 1, -11, -4, 69, -37, -73, 60, 75, -89, 4, 26, -95, 61, -15, 23, 60, -68, -8, 22, 22, 0, -64, 34, 77, 11, -87, -21, 110, -53, -61, -2, 62, 13, -6, 18, -3, -59, -30, 71, -37, -46, 78, -18, -11, 86, -87, -40, 17, -3, 73, 20, -2, 26, -36, -12, 36, -13, -35, 37, -66, 13, 10, -3, 51, -110, 40, 21, -56, -10, 73, 19, -59, 40, 20, -46, -6, 48, -1, 7, -42, -19, 47, -48, 7, 12, -59, 24, 86, 14, -48, -66, 26, 69, -68, -53, 74, 59, -30, -71, -42, 41, 36, 11, -29, -52, 77, 48, -3, -12, -32, -26, -32, -4, 15, 66, -14, -21, -1, -15, -4, 39, 5, 23, -3, -42, -8, -39, 19, 46, -17, -43, 91, 14, -8, -49, -15, 64, -2, 3, -59, -34, 65, -3, -36, -27, 62, 59, -49, -46, 42, 54, -11, -43, -10, -13, 4, 71, -76, 48, 3, -74, 27, -41, 76, -5, -90, 63, 36, 42, -71, 2, 6, -5, 0, -51, 78, 60, -83, -60, 13, 46, 82, 1, -83, -18, -14, 34, 29, -91, 85, 8, -29, -22, -6, 46, -53, 39, -25, 7, 80, -97, 11, 64, 8, 10, -76, -3, 69, -47, -86, 83, 22, -116, 86, 28, -44, 73, -48, 3, 3, -77, 15, 63, -9, 11, -2, -39, 49, -31, -7, -5, 5, 4, -54, 37, -8, -15, 14, 40, 47, -72, 12, 70, -56, -14, 9, -78, 37, 49, 17, 19, -3, -56, -7, 6, -68, 81, 57, -18, -39, -37, -24, 56, 56, -76, -17, 46, 18, -4, 0, -48, 55, 10, -91, 23, -23, 7, 35, 14, -30, -38, 32, 56, -3, 3, 63, -49, -5, 27, -48, -43, -31, 40, -8, 2, 76, -27, -40, 3, -31, 46, 69, -88, -51, 91, 21, -73, -7, 55, 48, -40, -71, -5, 10, 35, 0, -36, 6, -7, -26, 49, 37, -57, -18, 28, 57, 31, 22, -74, -55, 9, -25, -4, 12, 12, 65, 34, -39, -34, 0, 10, 13, 21, -18, 49, -56, 4, 9, -49, -3, -17, 2, 11, 38, -41, 62, 5, -96, 83, 17, -36, -36, -8, 69, -46, 31, 20, 8, -9, -13, 10, -1, 20, -82, 5, 45, -22, -10, 35, 39, -12, -93, 63, -3, -56, 48, -75, 62, 36, 9, -5, -113, 85, 74, -43, -53, 13, -2, -43, -14, 74, 56, -13, -17, -4, 12, -83, -26, 89, 65, -97, -36, 106, -58, -36, 52, -36, 23, -22, 26, 35, -53, 46, 6, -65, 2, 42, 39, -18, 0, 42, -36, -34, 47, -55, -37, 41, -47, 45, 20, -92, 58, 94, -97, -87, 58, 40, -10, -51, 44, 13, -18, 11, -51, -7, 35, 41, 35, -13, -70, 58, 2, 4, 23, -60, -23, -37, 72, 18, 11, -19, -52, 92, -58, -36, 90, 0, -81, -30, 60, 48, -18, -43, -49, 41, 36, -14, -7, -17, -32, 34, 18, -26, 42, 18, 28, -6, 2, 9, -76, 13, 77, -19, -6, -69, -30, 60, 21, -22, 29, -5, -64, 9, 38, -1, -58, -35, 95, 22, -75, 66, 56, -37, -53, 5, 1, -26, 0, 6, -40, 35, 20, -73, 19, 103, -52, -7, 49, -9, -11, -32, -12, 13, 68, 26, -97, 8, 100, -4, -58, -64, 81, -5, -99, 8, 93, -8, -14, -14, -1, 55, -2, 15, 3, -71, 2, 82, -81, -55, 77, -4, 0, 62, -80, -21, 87, -68, -14, 76, -49, -75, 14, 10, 10, 4, 21, -6, 18, 1, -24, 39, -56, -2, 32, 37, 36, -71, 9, 64, -15, -26, -29, 5, 11, 2, -13, -35, 68, -30, -68, 20, -17, 39, 11, -6, 66, -80, 8, 80, -80, 8, -15, 0, -20, 20, 36, 13, -26, -64, 79, 42, 21, -61, -39, 30, 49, -52, -113, 119, 3, -64, 8, -11, 82, 18, -106, 34, 46, 14, -17, -8, 19, -31, -9, 0, -10, 27, 12, -40, -13, -21, 26, -17, 7, 79, 17, -53, 23, 37, -45, -61, -28, 49, 37, -55, -40, 43, 66, 4, -30, -39, -3, 79, 17, -13, -10, -81, 12, 92, -32, 0, -39, -5, 94, -34, -15, 19, -66, 6, 37, -22, 35, 9, -59, -38, 64, -13, 7, 22, 13, -26, -20, 32, -60, 21, -3, 20, 28, 9, 21, -93, 8, 91, -99, -7, 57, -3, -8, -6, 2, 24, -5, -74, 36, 22, 1, -30, 32, 5, -10, 48, -21, -8, -32, -57, -7, 55, 52, 19, -23, -17, -53, -14, 51, -38, -42, 90, 69, -53, -5, -22, -4, -36, 18, 8, -11, 21, -21, 18, 25, -9, -44, 7, 69, 9, -49, -25, -26, 22, -28, 41, 95, -82, -60, 36, -10, 5, 14, -51, 63, 96, -69, -55, 81, -51, -45, 70, -52, 46, 65, -4, -56, -70, 23, -7, 31, 65, -57, 29, -25, -63, 71, 46, -32, 9, -28, -21, 14, -38, 61, -35, -28, -10, 23, 31, -60, -19, 77, 20, -88, 56, 18, -54, 76, 18, -37, 17, -7, -73, 23, 56, -24, -15, 12, -36, -27, 76, 29, -10, -46, -19, 65, 9, -28, -19, 42, 20, -40, 32, -74, 5, 64, -58, -25, 29, -38, 46, 24, -44, -24, 48, 9, -48, 35, 2, 25, 3, -9, -30, -8, 28, 60, -53, -45, 27, 34, -2, -62, 15, 4, -22, 2, 51, 32, -22, -31, 15, 22, -6, -29, -2, 43, -23, -28, -36, 5, -24, 57, 85, -55, -38, 23, 2, 14, -22, -78, 53, 60, -29, -37, -42, 57, 74, -103, 2, 48, -26, 15, -35, -28, 73, 73, -98, -36, 44, -45, 58, 20, -74, 29, 74, -1, -57, -12, 14, 8, 20, -43, -17, -10, 7, 31, 47, -29, -49, 47, 17, -49, -71, 93, 29, -108, 57, 41, -30, -30, 20, 26, -37, 80, -55, -51, 75, -2, -63, -20, 6, 46, 26, -28, 37, 53, -91, -3, 22, -29, 23, 21, 29, -48, 27, -54, -21, 60, -9, -53, 28, 10, -25, 13, -42, 31, 49, 36, -83, 7, 12, -74, 55, 14, 29, -20, -42, 75, -47, -17, 44, -27, 26, -38, -53, 31, 0, 17, 72, -8, -12, -14, 23, -40, -22, 95, -10, -60, 13, 40, -74, 7, 78, -19, -63, -4, 70, 6, -65, 44, -11, -19, 19, -8, 53, -35, -87, 55, 93, -18, -42, -10, -9, -41, 38, 77, -60, -58, 18, 44, 70, -55, -37, 57, -76, 10, 30, -5, 17, -31, 38, 2, -28, -57, 15, 4, -1, 41, -53, 4, 21, 14, -25, -10, 86, 10, -22, -63, -51, 106, -20, -91, 53, 31, 56, -22, -47, -1, -26, 55, 78, -100, -30, 48, -44, -35, 31, 70, -19, 3, -39, 23, 15, -68, 36, -12, -34, -6, 14, 4, 79, -5, -62, 20, 47, -10, -1, 1, -12, -7, -56, 68, -20, 28, -14, -63, 102, 14, -83, -5, 15, -10, 0, 11, 32, 12, 3, 0, 1, 37, -87, -6, 29, -41, 14, -55, 85, -10, -53, 73, -42, 28, 4, -39, 54, -11, -81, 45, 3, -53, 19, 0, 49, -6, 35, -6, -86, 59, -34, 32, 75, -119, 28, 79, -23, -92, 49, 56, -104, 21, -6, -9, 28, -22, 63, 60, -32, 5, -8, -7, -48, 10, -7, -2, 24, -83, -5, 29, 63, -40, -24, 24, -26, 3, -25, 61, -1, 27, 6, -83, 48, -22, 19, 53, -21, -7, 20, -36, -3, 14, -66, 61, 2, -72, 63, 5, -42, 34, 38, 19, 12, -75, -65, 97, 12, -89, 48, 34, -63, 32, 63, -15, -80, -4, 32, 5, -9, -76, 83, 74, -83, 41, 23, -60, -7, -48, 58, 37, -14, 8, -31, -2, 18, 13, -35, 31, 56, -96, -42, 103, 44, -89, -22, 76, -6, 12, -25, -18, 66, -57, -30, 4, -14, -29, 35, 66, -77, 7, -10, 40, -6, -42, 36, 10, -26, 2, 45, 7, 15, 0, 20, -31, -65, -2, 22, 42, -12, -4, 44, -57, -37, -8, 39, 36, -39, -12, -8, -5, 83, -18, -54, -36, 52, 71, -25, -64, -17, 19, 53, 0, -90, 75, 55, -44, -37, -9, -6, 61, -14, -71, 5, 37, 8, 46, -36, -6, 31, -49, 9, -15, 47, 42, -54, 8, 24, -81, 53, -12, -59, 109, -39, -17, 72, -73, -41, 11, 7, 65, -58, -3, 104, -55, -55, 22, -11, 20, -6, 23, -27, 1, 26, -95, 48, 60, 26, -60, 4, 78, -78, -30, 51, 18, -47, -9, 59, 0, 1, -23, -25, -36, -29, 58, 0, 6, 58, 11, -63, -38, 31, 18, -57, 40, 35, -11, 12, -28, -53, 20, 24, -19, -7, -35, 0, 31, 64, -52, -53, 65, 11, 12, 7, 6, -20, -85, 35, 15, 19, 60, -22, -34, -35, 55, -17, 0, 43, -3, -27, -9, 15, -3, -27, -12, 71, -29, -69, 24, 27, -9, -41, 63, 0, -32, 73, -46, 19, -26, -9, 58, -79, -6, -2, 0, 25, -19, 0, 69, -21, -27, 58, -4, -31, 28, 3, -72, 0, 24, 41, 28, -75, -90, 94, 9, -8, 32, -11, 6, 4, 4, -70, 37, 86, -71, -51, 0, 20, 62, -66, 23, 31, -7, 19, -2, 41, -91, -51, 18, 45, -5, -83, 82, -7, 13, -18, 3, 43, -31, 35, -64, -27, 75, -27, -52, 5, 12, 37, 28, -37, -8, 52, -5, 3, -44, 17, 22, -21, -56, 42, 25, -87, 96, -26, -71, 107, -46, -41, 14, 35, 80, -48, -77, 42, 35, -42, 51, -63, 15, 77, -103, 32, -7, 26, 13, -51, 43, 36, -74, -10, 81, -72, 37, 41, -74, -10, 11, -7, 36, 26, -61, 25, -25, -26, 46, 10, -45, -39, 83, -51, 18, 93, -19, -81, 29, -7, -20, 54, 6, 41, -74, -1, -9, -36, 20, 6, 45, 8, 20, -9, -56, -17, -5, 10, 43, 43, -90, 20, 3, -29, 82, 18, -26, -26, -40, -19, 54, 51, -78, -24, 90, -40, -45, 58, 36, -28, -23, -8, 0, -2, -39, 36, 68, -45, -41, 22, -5, -21, 22, -1, -28, -5, 17, 32, 57, -21, -76, 21, 27, -45, 0, -14, 27, 62, -68, -21, 32, -2, 58, 35, -95, -72, 72, 63, -27, 30, -25, -9, 7, -3, -13, -19, -6, 1, 34, -62, -17, 48, 52, -13, 30, -63, -7, 59, -26, 59, -77, -79, 54, 90, -65, -37, 17, 5, 26, -8, 35, -2, 1, -68, -1, 77, 0, -8, -7, -75, 39, 61, -25, 1, -40, 2, 45, -48, -48, 44, -11, -36, 54, 45, -56, 9, 5, -38, 13, 30, -47, 51, 30, -47, -17, 29, 28, -15, 24, -3, 41, -48, -31, 38, -74, 42, 19, -25, -3, -31, 19, -38, 47, 53, 6, 8, -29, -75, -29, 74, 45, -74, 14, 77, -12, -4, 18, -75, 0, 40, -75, 20, 78, 7, -74, 29, 48, -54, 5, 21, 24, 23, -106, -18, 72, 11, -4, -90, 48, 54, -12, -15, -1, 21, -53, 9, 17, -57, 47, -4, -35, 86, 13, -46, 0, -41, -14, 27, 13, -9, -63, 63, -10, -56, 27, 40, 68, 0, -25, 24, -39, -18, 6, -38, -17, 45, 62, -23, 13, -3, -7, -2, -32, 26, -47, -52, 75, 24, -22, -17, 12, 47, -88, 3, 99, -60, -44, 75, -41, -71, 80, 7, 24, -45, -4, 2, 1, 58, -23, 36, -60, -7, 9, 21, -4, -38, -5, -39, -11, 60, 32, 1, -4, -32, 26, -39, 18, 93, -96, 1, 19, -17, 31, -93, 75, 2, -88, 78, 35, 25, -22, 0, 15, -11, 21, 12, -52, 12, -24, -64, 74, 5, -41, -42, -23, 77, 5, -3, 59, -68, -6, 79, -82, 4, 100, -32, 28, -79, -47, 85, -55, -66, 64, 51, 31, -26, -25, 3, -35, 37, 49, -72, -42, 8, -24, 24, 62, 4, -68, 10, 44, 36, -44, -14, 61, -57, -22, 64, -24, -66, 14, 32, -23, -34, -2, 9, 28, 63, -9, 15, 8, -48, -55, 56, 49, -82, -5, 2, 31, 13, 11, -12, -40, -11, -26, -1, 22, 42, 41, 0, -4, -30, -79, 85, 21, -81, -17, 74, -20, -25, 91, -10, -76, 35, 46, -26, -44, 20, 87, -17, -56, 11, -28, -8, 93, -78, 13, 2, -14, 54, 0, 3, -90, -55, 64, 22, -45, 51, -14, -43, 22, 54, 56, -56, 1, 13, -87, 63, 36, -108, 48, 69, -6, 19, -28, -4, -41, -17, -2, -55, 40, -22, 39, 38, -76, -3, 61, -11, 23, 48, -36, -44, 12, 17, 10, -6, 10, 60, -57, -42, -27, -11, 25, -30, -12, 89, 54, -51, -37, 51, 4, -22, 49, -43, -94, 83, 37, -30, -17, -25, 15, 31, 41, -81, -36, 48, 21, -25, 0, -32, 19, 62, -62, 47, 28, -54, 44, -10, -87, 9, 17, 28, -8, -66, 96, 5, -92, 26, 87, -23, 0, 14, -81, 41, 19, -7, -18, -68, 77, 69, -100, 9, 19, -29, 34, 46, -63, -31, 40, -62, 68, 36, -28, 57, -9, -20, -51, 29, 2, -78, 31, -18, 26, 38, 22, -42, -57, 3, 0, 0, 51, 12, 10, -41, 3, 43, -15, 52, 9, -87, 13, 76, -53, 5, 17, -36, -39, 79, -29, -34, 4, -20, 58, 30, -68, -30, 98, -38, -24, -10, -15, 24, 0, -6, -15, 6, 35, -10, -54, 45, 11, -38, -10, 70, 78, -105, -57, 61, -48, 26, 3, -40, 6, 61, -9, -63, 57, -47, 32, 8, -58, 18, 10, 58, -13, 15, -27, -69, 7, 7, 68, -3, -7, -32, -22, 68, -46, 12, 107, -74, -49, 0, -3, 46, 43, -15, 4, -11, -42, 38, -24, 13, 29, 8, -19, -73, 24, 41, -49, 13, 51, 14, 34, -71, 2, 11, -26, 88, -90, -6, 14, -48, 81, 11, -93, 35, -4, 23, 0, -43, 60, -27, -7, -20, -18, 63, -3, 8, -7, -35, 43, -70, 6, 52, -26, -11, 61, -30, -36, -2, -61, 72, 37, 22, -28, -32, 55, -32, -8, 55, -56, -61, 28, 25, 7, 11, -22, 27, 19, -29, -3, 41, 11, 0, 2, -106, 10, 42, -46, 66, 18, -82, 23, 77, -61, -3, 44, -8, -14, -78, 48, 19, -45, 58, 43, -17, -21, -69, 11, 86, 11, -104, 37, 43, -103, 20, 27, 0, 42, 4, -21, -54, 52, 1, -85, -6, 88, 47, -10, -40, -7, 35, -24, -31, -17, 23, 39, 48, -45, -38, 46, -36, -31, 63, -13, 3, -52, 39, 2, -9, 41, -21, -38, -38, 94, -37, -43, 71, 29, -36, -79, 23, 87, -11, -7, -20, -81, 54, 4, -12, -5, 31, 62, -39, 6, -41, -39, 68, -24, -35, 58, 17, -57, 18, -19, 15, 93, -65, 0, 9, 7, 30, -78, 7, 15, 23, -32, -62, 78, -51, 37, 71, -109, 9, 30, -11, 59, -5, -56, 54, -21, -111, 73, 11, -2, 53, -60, 0, -15, 51, 8, -117, 83, 15, 2, -8, -66, 80, 17, -8, 51, -38, -31, -32, -48, 88, 65, -104, -6, 34, -73, 62, 14, -22, 96, -80, -58, 36, 4, 39, -45, 14, 55, -76, -54, 55, 1, -6, 1, 41, 1, -57, 6, 58, -1, -44, 59, -48, -11, 28, -38, 51, -42, 0, 51, -81, 31, 79, -46, -47, 7, 19, 56, 39, -34, -87, -15, 79, -7, -12, 10, -4, 39, 13, -35, -53, -5, 0, -10, 73, 8, -23, 9, -11, -24, 34, 40, -103, 5, 106, -64, 11, 35, -98, 74, -23, -71, 37, 36, 31, 22, -40, -64, 85, -49, 11, 7, -54, 14, -2, 18, 23, -25, 26, 11, -49, 63, 26, -19, -41, 20, 48, -30, -56, -24, 20, 13, -8, 57, -37, -64, 78, 8, -12, 27, -18, -1, 35, -72, 12, 32, -55, 37, 7, -27, 45, -19, -74, 75, 48, -4, -15, 8, -15, -75, -14, -15, 30, 69, 19, 15, -86, 4, 43, -103, 35, 4, 9, 49, -64, 23, 58, 14, -53, -21, 8, -28, 47, 45, -66, 9, 61, -87, 20, 21, -45, -18, 7, -13, 49, 26, 0, -11, -78, 44, -26, 45, 49, -105, -14, 95, 27, -68, 21, -26, 22, 8, -58, 96, -80, 10, 79, -19, -52, -12, 5, -7, 61, -8, 0, 21, -72, -1, 96, -39, -66, -19, 6, 74, -36, -5, 58, 11, -54, -31, 8, -56, 65, 65, -93, 9, 72, -13, -7, 21, -26, -3, 35, -80, 9, 12, 31, 49, -102, 39, 7, -54, -1, 14, 21, -38, 31, -34, -24, 68, 25, -38, 35, 1, -88, 75, -11, -10, 60, -22, 31, -81, -2, 42, -46, -13, 55, 5, -76, -20, 22, 22, 15, 1, 41, 34, -14, -38, 19, -19, -83, 44, 55, -70, 25, 79, 4, -75, -22, 62, 12, -11, -13, 10, 29, -61, -3, 83, -56, -77, 42, 77, -57, -29, -13, 5, 4, -52, 78, 3, -90, 109, 25, -36, 58, -39, -44, 58, -6, -64, 12, 5, 30, -2, -91, 62, 42, -92, 14, 99, -60, -51, 70, -5, 5, 35, 1, 6, 7, -34, 31, -64, -37, 57, 11, 0, 15, -9, -51, 8, 35, -61, 17, 71, -89, 61, -2, -41, 78, 8, -29, -73, -22, 14, 34, -15, -60, 37, 78, 59, -107, 22, -6, -34, 56, 5, -9, -38, -1, 25, 81, -99, -9, 96, -31, -74, 24, 76, -5, -7, -2, -39, 31, -45, -23, 66, -83, 29, 102, -95, -2, 17, -95, 81, 74, -39, -1, -27, -59, -3, 0, 0, 8, -7, -35, 92, 5, -10, 78, -92, 2, 52, -15, 9, 4, -11, -59, 55, 14, -69, -15, -8, 37, 0, -34, 0, 73, 53, -47, 14, 47, -25, -75, -56, 78, -20, 12, 107, -126, 3, 12, -10, 31, -2, 21, -74, -14, 74, -38, -21, 119, -78, -4, 43, -78, 68, 42, -95, 28, 15, -81, 56, 82, -65, 3, 49, -69, 38, 19, -56, 15, 31, -44, -62, 31, 65, -47, 20, 27, -68, 21, 9, -9, -7, 32, 45, -54, -13, -27, -47, 96, -18, 9, 66, -64, 34, 2, -110, 72, 0, -52, 68, 11, 15, 3, -44, -10, -25, -25, 0, -1, 86, -11, 11, -13, -68, 57, 19, 11, 7, -3, -7, 9, 26, -55, -29, 38, 35, -24, -23, 56, -57, -69, 91, -44, -62, 26, 37, 3, -20, 37, 22, -26, -63, 32, 47, -20, -20, -20, 10, -14, -25, 4, -22, 94, 36, -54, 45, -20, -61, 23, 17, -28, 69, -26, -48, 3, 1, -8, -15, 93, 25, -80, -45, 73, 41, 2, -36, -70, -19, 63, 7, -63, 66, 2, -56, -7, 60, 76, -28, -86, -13, 97, -5, -54, -37, 56, 37, -57, 46, 42, -54, -40, 71, 11, -78, 22, 15, -25, 41, -1, -73, 48, 45, -5, -57, -10, 95, 0, -22, -47, 44, -36, -60, 40, -3, 17, -35, 34, 92, -105, -10, 37, -30, 39, 26, 22, -52, -46, 19, -30, 39, 58, -94, -1, 49, -41, -12, 30, -13, -59, 98, 5, -94, 42, 24, 14, 32, 9, -39, 12, 37, -52, -61, 26, -13, -30, 30, 22, 11, 29, 13, -38, -24, 30, 49, 3, 12, -55, -53, -5, -3, 24, -18, 18, 41, 27, -57, -13, 34, 12, 0, -37, -38, 26, 82, -75, 20, 0, -28, 26, 29, -13, -14, 28, -95, 58, 29, -81, -17, 69, 1, -15, -17, 4, 0, 23, 30, -57, 9, 63, -19, -103, 28, 29, 37, -21, -21, 53, -22, -27, -31, 7, 72, -64, 13, 86, -5, -65, 27, -25, 2, 28, -41, -11, 9, 71, 8, -46, -77, 40, -4, -6, 28, 2, 47, -47, 4, 25, 4, -19, -1, -26, -11, 70, -93, 27, 21, 10, 73, -85, 10, 74, -57, -31, 59, -23, -73, 71, 17, -36, -24, 37, -44, 5, 38, 0, -19, -69, 27, 72, 23, -86, -39, 9, 72, -41, 15, 117, -123, 0, 28, 0, 51, -28, -7, -1, -53, 29, 47, -32, -6, 25, 2, -49, 31, 40, -49, 12, -28, -21, 87, -27, 7, 21, 8, -34, -1, 46, -54, 11, 20, -23, 35, -42, -30, 26, -65, 31, 34, -14, -1, 28, 8, -3, 1, -72, 38, 64, -81, 9, 63, -109, 7, 44, 24, 17, -102, 48, 38, -43, 62, -52, -42, 72, 17, -70, -32, 64, 46, 3, -40, -46, 54, -35, -47, 32, 4, -6, -37, 59, -17, 6, 61, -11, -37, -2, 2, -24, 21, 41, -44, -29, -9, 24, 23, -12, 64, -9, -37, 18, 12, -79, -24, 44, -22, 19, 57, -13, 10, 39, -46, -99, 68, -9, 4, 9, -11, 8, -14, 10, 27, 49, -18, -72, -15, 2, 26, 27, -7, 9, -65, 7, 20, 1, 29, 19, -70, 0, 1, 52, 17, -43, -20, -48, 59, 70, -39, -39, -31, 55, 80, -119, 20, 58, -78, -14, 41, 61, 9, -54, -40, 56, 40, -20, -31, -17, 0, -13, 70, 3, -49, -3, -41, 18, 39, 19, -23, 23, -23, -55, 81, 29, -38, -10, -19, -3, 60, 22, -32, -19, -35, 36, 38, -105, 18, 93, -9, -93, -7, 57, 21, -56, -77, 93, 49, -38, 22, -60, -15, 86, -4, -46, 26, -22, -57, -13, 83, 2, -100, 54, 71, -24, -18, -3, 1, -2, -18, -4, -5, 62, 53, -94, 6, 87, -4, -31, -40, 13, 17, -58, -8, 12, 5, 0, -29, 60, -14, -54, 64, -8, -1, 24, -11, -21, 21, -9, -24, 3, -36, 80, 65, -93, 6, 70, -8, 23, -75, -26, 18, 34, 5, -13, 70, -102, 8, 38, -40, -6, -17, 22, -14, -14, 24, 85, -41, -41, -35, 44, 48, -71, 36, 1, -32, 41, -40, -18, 43, -23, 44, 60, -79, -41, 70, -34, -27, 57, 5, -70, 49, -9, -47, 36, -27, 0, -12, 44, 45, -48, 0, -17, 13, 11, -13, -15, 32, 57, -39, -12, -57, 27, 23, -26, -11, -36, 54, 45, 22, -51, -2, 70, -62, -26, -27, 21, 60, -39, -20, -5, 23, 68, -24, -51, -9, -41, 43, 0, 19, 6, -36, 76, 9, 10, -60, 0, 82, -9, -43, 13, -40, -46, 63, -12, 15, 37, -79, -11, -1, -11, 70, 21, -35, -42, -29, 44, 8, -7, 45, 26, 21, -83, 9, 51, -74, -51, 51, -13, 52, 8, -109, 12, 48, 43, 1, -20, -29, 31, 53, -31, -69, 35, -9, -14, 81, -40, -59, -20, 62, 95, -107, -2, 9, 15, 24, -63, -30, 53, 59, -113, 62, 58, -103, 26, -7, 9, 95, -39, -45, 37, 38, -5, -40, -61, 0, 18, -7, 30, -1, -31, 13, 4, 51, 22, -65, -35, 69, 11, -90, 14, 32, -46, 52, 41, -21, -46, -39, 73, 1, 27, -1, -48, 22, 45, 1, -89, -22, -7, 32, 64, -40, -42, -20, 10, 69, 3, -20, 27, 13, 21, -69, -66, 109, -40, -22, 88, -90, -37, 23, 48, -32, 23, 0, -9, 72, -23, 38, -88, -4, 66, -23, -41, 0, 69, -32, -20, -19, -32, 6, -26, 81, 25, -90, 78, 3, -90, 32, 28, -38, 36, 77, -49, -31, -13, -37, 12, 78, -22, -73, 77, 20, 14, 32, -66, -5, 0, 1, 63, -29, -104, 60, 49, -79, -4, -5, 40, -6, 5, 70, -23, -46, 32, 55, -81, -89, 20, 20, 80, -24, -26, 44, 15, 8, -37, -27, -20, 75, -24, -66, 44, -14, -26, 74, 15, -34, -17, -58, 89, -13, -97, 65, 48, -61, -8, 80, -64, 10, 14, -95, 98, 75, -51, 25, -6, -66, -25, 85, -14, -47, 21, 8, 47, -8, -5, -25, -43, 61, 29, -61, -61, 42, 94, -35, 3, -6, -46, -39, -17, 57, -22, -26, 21, 58, -27, 17, -7, -54, 104, -24, -79, 10, -17, 81, -17, -21, 54, -63, 65, -49, -10, 91, -7, -5, -35, 19, -36, 8, 69, -51, -41, 46, 29, -23, 17, -87, -5, 94, -28, -11, -39, 3, 86, -53, -26, 87, -56, -86, 47, -15, -21, 13, 75, -6, -106, 42, 99, -28, -57, 56, 52, -102, -5, 81, -12, -11, -5, 2, -31, -8, -35, 40, -2, -81, 97, 80, -102, -70, 105, 32, -82, -28, 69, -6, -57, 75, 31, -45, -45, -4, 10, -18, 7, -15, 64, -5, -28, 60, -1, -59, 28, 76, -20, -88, 18, 77, -27, 27, 4, -13, -30, -79, 70, 14, -85, 35, -20, -49, 79, 23, -55, -18, 7, 63, -37, -36, 59, 41, 23, -53, 3, 72, -89, -15, 94, -72, -49, 88, -45, -40, 54, 10, -6, -6, 30, 19, 4, 10, -9, -6, -55, -64, 61, 43, -20, 23, 28, -53, -23, 51, 2, -21, 10, -63, -36, 85, -46, 27, 38, -71, 9, -39, 54, 89, -47, -3, 17, -22, 3, 7, -51, 39, 55, -102, -3, 52, -77, 4, 89, 11, -57, 1, 12, -69, 27, 70, -4, 4, 4, -57, -44, -10, 15, -10, 58, 80, -19, -12, -32, 6, -29, 26, 47, -87, -48, 19, 58, -36, 26, 37, -4, -10, -73, 12, 5, 66, -28, -87, 72, 65, -52, 5, 58, -39, 14, 26, -52, 13, 10, -81, 1, 93, -57, -59, 9, -15, 52, 45, -31, -12, -4, -36, 63, 9, -23, -17, -34, 60, -14, 38, 12, -48, 65, -40, -68, 79, -36, -3, 73, -24, -64, -38, 72, -31, -8, 60, -26, -45, -3, 52, 28, -32, 43, -20, -1, 17, -38, -9, -60, 81, 3, -44, 58, -65, 26, 79, -7, 13, -15, -25, -8, 7, 48, -72, -1, 39, -9, -28, -7, -14, 25, 23, -47, 68, 0, -25, -28, -36, 51, 22, -64, -32, -24, 82, -6, 3, 72, -109, 40, 32, -22, 29, -70, 25, 69, -71, -43, 57, 11, -72, 44, 36, -53, 20, -9, -27, -27, 52, 24, 24, -31, -40, 102, -56, -69, 94, 56, 2, -104, 6, 31, -14, 15, -37, 36, -51, 4, 78, 9, -94, 27, 54, -57, -23, 52, 46, -77, 47, -12, -28, 71, -48, -45, 37, 6, -4, 20, -23, -5, 27, -38, 28, 11, -23, -6, 25, 60, -116, 14, 69, -100, 44, -11, -20, -1, 40, 24, -77, 90, 9, -83, 25, 72, -20, -46, -8, -4, -51, 61, 80, -23, -66, 18, -11, 20, 11, -98, 79, 5, -78, 18, 18, 56, -13, -3, 75, -64, -69, 17, 2, 29, 45, -82, 17, 23, -19, -11, -2, 62, -65, -9, 37, -21, -12, 27, 0, -23, 44, 59, -18, -12, -37, 22, 40, -54, 45, -21, 15, -47, -1, 18, -18, 44, -63, 0, 44, 28, -12, -45, -20, 31, 35, -1, 9, 40, -65, -76, 12, 86, -18, -114, 74, 53, -91, 5, 0, 39, 98, -115, 14, 94, -97, 21, 1, -28, 21, -61, 0, 98, -17, -20, 42, -75, -2, 54, -56, 22, 66, -38, 0, 45, -22, -37, -9, -1, 55, -11, -48, 41, 3, -32, 1, 40, -34, 5, 12, -31, 54, 10, -22, -55, 14, -5, -17, -7, 26, 40, 13, 3, -90, 36, 23, 0, -22, 11, 20, -76, 2, 61, 53, 6, -59, -36, 43, 17, -28, -55, 4, 24, -39, -37, 59, 62, -39, -68, 77, -15, -26, 93, -36, 15, 15, -100, 17, 80, 23, -72, -83, 22, 97, -28, -79, 39, 44, -36, -54, 15, 0, 43, 19, -39, 28, -30, 21, 97, -98, -8, 79, 4, -29, -46, 44, -39, -34, 39, 44, -6, -56, 73, 13, -45, -69, 45, 82, -42, 12, 26, -7, -81, -17, 13, -30, 99, -19, -95, 86, -9, 6, 53, -94, -1, -17, 43, 49, -52, -5, -15, 49, 46, -53, -24, 0, -13, 20, -26, -34, 31, -21, 52, 41, -38, -46, 34, 57, -66, -35, 5, 59, -52, 38, 78, -56, -66, 32, -5, -30, 115, -22, -66, 52, 30, 15, -58, -69, 37, 2, -12, 47, 3, -49, -21, 75, 12, -98, 24, 56, -45, 32, 2, -75, 74, 59, -20, 5, -20, -6, -4, -14, -30, 37, 38, -110, 58, 66, -69, -13, -42, 54, 8, -35, 3, -13, 42, -7, 23, -44, -62, 89, 76, -60, -77, 61, -1, 12, 44, -20, 28, -74, -14, -3, -32, 0, 1, 4, 45, 46, -35, 29, -11, -4, -9, -8, -18, 34, -13, -18, 102, -78, -15, 64, -27, 18, -6, -8, 52, -75, -6, 56, -36, -41, 32, 42, -63, 34, 69, -110, -7, 29, 27, -19, -86, 21, 60, 10, -79, 69, 10, -89, -7, 83, 68, -36, 11, -32, -23, 39, 2, -28, -12, -34, 41, -1, 9, -1, -79, 81, -24, 24, 0, -105, 119, 2, -80, 68, 9, -24, 3, 23, -4, -7, 17, -28, -22, 4, 51, -45, -64, 55, 14, 10, 24, -54, 29, 31, -56, -24, -22, 36, 90, -45, -43, 94, -22, -102, 27, 98, -18, -80, 36, -24, 20, 30, -49, -1, 37, 0, -45, -25, 31, 81, -17, -31, -63, 13, 89, -30, -6, -45, 25, 80, -93, 5, 41, -2, 11, -42, 8, -6, -12, 21, -28, 11, 29, 30, 9, -21, -59, -37, 41, 63, 41, -65, -57, -23, 62, 7, -52, 54, -40, -1, 0, 4, -21, 42, 1, -7, 3, -12, 94, -9, -80, -24, 1, 59, 5, -99, 40, 34, -25, -29, 9, 17, -4, 41, -4, -54, 49, 55, -23, 32, -59, 0, 32, -80, 42, 32, -89, 46, 22, 4, 35, -57, -18, 36, 4, -35, 49, 19, 25, -90, 10, 34, -73, 6, 54, 35, -48, 12, 0, -51, 19, 54, -48, -78, 88, 82, -65, 22, 14, -23, 47, -62, -58, 27, -47, 37, 83, 2, -31, -5, 44, -22, -80, -28, 96, -49, 9, 46, -37, 11, -6, 4, -70, 59, 36, -94, 54, -9, -71, 45, 80, -46, -13, 25, -42, 71, -52, -44, 71, 24, -49, 6, 4, -43, 93, -34, -68, 103, 8, -83, 1, 4, 8, 43, -45, -64, 62, 97, -97, 11, 52, -108, -12, 13, 9, 37, 62, -20, -98, 45, 2, -37, 30, -14, 57, -10, -27, 8, -21, -15, 13, 69, -11, -63, 2, 51, -19, -44, 36, 18, -54, 66, 22, -66, -26, 30, 100, -77, -97, 114, 55, -93, -34, 85, 23, -90, -13, -5, 7, 55, -44, 47, 11, -34, -19, 13, 21, -59, 81, 32, -18, -64, 11, 3, -43, 73, 38, -51, -6, 72, -52, -40, -22, 27, 23, -21, 51, -14, -3, -28, -74, 86, -4, -61, 54, -46, 65, 51, -83, 57, -5, -102, 80, 93, -95, -51, 75, -59, 10, 46, 11, -40, 6, -9, -13, 28, -30, 38, 14, -31, -15, 76, -82, 3, 15, -53, 92, -55, 22, 7, 2, 15, -97, 108, -25, -58, 35, 28, 14, -69, -10, 26, 1, -27, 19, -10, 2, -11, 27, 18, -46, 35, -41, 7, 14, -46, 69, 83, -78, 0, 0, -75, 103, 14, -77, -34, 71, 44, -2, -24, -2, -17, 2, 0, -43, 23, -34, 73, -12, 15, -22, -37, 48, -64, -25, 43, 0, 41, 13, -55, 41, -8, 3, 8, 8, 36, -26, -8, -9, -10, -34, -34, 63, 59, -34, -68, -29, 42, 93, -38, -51, 70, 37, -23, 4, 28, -74, -83, 72, 28, -24, -22, 44, -21, -12, 52, 12, -17, -69, 3, 61, -11, -31, 38, -64, 46, 59, -96, 1, 37, -2, -52, -1, 34, 31, 3, -44, -39, 31, 2, -9, 8, -19, 34, -13, -9, -23, 0, 62, -2, 4, 12, 5, -3, -85, 75, 17, -22, -19, 19, 17, -45, 77, 14, -99, 19, 19, -56, 71, 29, -26, -49, 37, 61, -15, -63, -60, 72, 22, 2, -21, -63, 38, -37, 22, 64, -74, -46, 41, -4, 62, 37, -25, 49, -63, 6, 47, -42, -27, 5, -10, 31, 69, -85, 4, 48, -37, -54, 8, 8, -73, 80, 36, -59, 65, -28, -107, 102, 9, -64, 11, -38, 80, 93, -98, -68, 99, 36, 1, -41, -47, 9, -9, 0, 38, -4, -60, 2, 30, 40, -11, -18, 7, 44, -56, -60, 127, -53, -68, 27, -5, 29, -10, -10, 9, 0, 30, -2, -52, 31, 46, -8, 41, -54, -99, 81, 30, -69, 63, 62, -6, -41, -49, 22, -19, -13, 76, -27, -41, 8, -22, 64, 12, -7, -59, 45, -11, -27, 43, -63, 4, 64, 62, -65, -79, -15, -6, 42, 4, 56, 14, -91, 13, 56, 21, -5, -45, -13, 79, 0, -4, -32, -27, 30, -66, 25, 55, -75, 0, 75, -25, 3, 48, -54, -61, 60, 17, -64, -7, 44, -8, -14, 65, 2, -48, -2, -3, 14, -15, -34, 14, 68, 23, -9, -12, -21, 15, 17, 37, -98, 5, 8, 15, 34, -47, -19, -39, 83, 2, -46, 17, 13, -42, -28, 19, 0, 60, -5, 15, 42, -18, -62, 17, 24, -74, 6, -19, 56, 4, -1, 69, 7, -83, -2, 39, -17, -44, 1, 66, -46, -19, -48, 81, 25, -77, -8, 25, 94, -17, -48, 45, -37, 1, 40, -10, -70, 25, 81, -17, -60, -11, 76, -76, 18, 48, -35, 1, 1, -10, -43, -41, 58, -1, 19, 83, -57, -81, 19, 32, 9, -26, -52, 86, 61, -8, -36, 10, 37, -69, 14, -23, -78, 66, 10, -55, -13, 90, 31, -11, -28, -11, 55, 5, 8, -17, 1, -51, 11, 0, -15, 24, -53, 68, -2, -80, 57, 71, -70, -19, 26, -76, 47, 41, -27, 60, -18, -23, 59, -78, -11, 5, 20, 43, -100, 55, 1, 10, 4, -95, 10, 80, 19, -39, 37, 12, 12, -21, -5, -37, -39, 0, 0, -12, 17, 107, -64, -90, 105, -29, -55, 69, -24, -7, -22, 10, 20, -18, 24, 3, -1, 34, -6, -74, 17, 3, 53, 7, -12, 48, -30, -53, 27, 82, -70, -19, -34, -23, 91, 25, -27, -52, -17, 58, 24, -35, -38, 44, 55, -17, -41, -36, 15, 40, 2, -79, -43, 53, 39, -57, -6, 7, -1, 23, -39, 43, 91, -76, -65, 72, 59, 15, -92, -45, 74, 20, 30, -76, -22, 83, 14, -62, -60, 34, 64, 29, -42, -64, -27, 106, -36, -30, 5, -36, 102, -38, -80, 83, -5, -38, 44, -31, -24, 37, 37, -61, -29, 65, -28, -51, 40, -10, -23, 69, 20, -45, 10, -21, -25, 97, -48, -37, 68, -70, 61, 35, -83, 1, -15, 26, 52, 4, 17, -63, -46, 53, -36, 14, 100, -65, -12, 27, -78, 74, 73, -35, -60, -27, 53, 25, -64, 28, -12, -20, 94, -64, -74, 8, 26, 0, 37, -32, 25, 52, -95, -19, 85, -20, -4, 74, -66, 4, -35, -7, 56, 40, -42, -8, 34, -102, 20, 61, 14, 7, -45, -2, 54, -32, 8, -30, -10, 44, -63, 14, 74, -47, -2, 48, -48, 13, -13, 21, -5, -46, 12, 51, -4, -30, 44, 5, 1, -48, -22, 39, -63, 46, 12, -11, 36, -91, -18, 2, 46, 8, 19, 9, -19, 35, -55, -43, 25, 43, -44, 22, -2, -31, 73, -9, -40, 5, 19, -61, 48, 90, -44, 6, 21, -9, 19, -76, 11, 89, -75, -31, 8, -55, 66, 79, -19, -79, -55, 6, 55, -6, 8, 52, -19, -6, -68, 51, 85, -47, -100, 43, 41, -35, 51, -51, -22, 46, -14, -7, 2, 48, -64, -9, 107, 0, -20, -1, -78, 13, 92, -23, -81, 13, 26, 9, -13, -42, 83, -41, -91, 96, -19, -48, 61, 7, 34, -74, -30, 20, 2, 83, -63, -38, 94, -73, -12, 53, 12, 18, -44, 20, -6, -14, 10, 21, -4, -5, 3, -54, 63, 23, -93, 71, -27, -31, 81, -19, 28, -64, -87, 32, 108, -62, -2, 91, -116, 5, 6, 35, 0, -36, 55, -7, -27, -46, 13, 58, 37, 17, -86, 11, 38, -68, 62, 8, -76, 28, 13, -70, 55, 18, -35, 52, -23, -15, 5, 0, -35, 14, 32, -37, 4, -46, 66, 63, -93, -6, 28, -32, -13, 57, -40, 3, 102, 18, -75, -64, 46, 26, -20, -29, 45, 76, -93, -64, 60, 3, 22, 25, -69, -56, 99, 21, -100, 59, 85, -61, -60, 2, 17, 15, 37, 0, -71, 48, 13, -35, -37, 63, -7, -58, 34, 37, 15, -58, -25, 53, 58, -3, -32, 10, -41, -45, 32, -30, 15, -15, 20, 46, -35, 59, -30, -86, 56, 9, -57, 51, 87, -97, 7, 75, -25, -70, 4, 100, -40, -19, 64, -74, -2, 30, -83, 46, 75, -48, -72, -19, 45, 37, 3, 36, -15, -6, -30, -71, 4, -1, 73, 72, -76, -10, 37, 6, 28, -70, 18, 7, -93, 64, 24, 18, -37, -35, 63, 17, 29, -32, 19, -15, -87, 45, -4, 10, 18, -55, 54, -1, -32, 36, -44, 25, 1, -8, 56, -83, -54, 53, 12, -30, -13, 39, 95, -53, -83, 66, -17, -56, 36, -19, 19, 43, 3, 37, -37, -70, 3, -5, 20, 64, 8, -1, -23, 31, 11, -104, 63, 43, -47, -31, 10, 46, 6, -5, 14, -54, -75, 112, -22, -56, 95, -5, 6, 6, -57, -30, 24, 37, -36, -44, -8, 87, 41, -34, 30, -60, -4, 70, -13, -30, -78, 19, -6, 43, -5, -12, 100, -79, -11, 76, -3, -30, -19, 24, -45, 15, 83, -22, -31, -63, 41, 66, -89, -5, 54, -82, 48, 26, -9, 36, -26, 46, -80, -8, 88, -89, 0, 52, -31, -12, 14, -12, -46, 0, -10, 17, 14, -35, -1, 69, 12, -69, 26, 31, 36, -51, -24, 82, -26, -12, 3, -28, 8, 36, -37, -35, 60, 73, -95, -58, 60, 8, 19, -6, 11, 9, 11, 23, -6, -82, 4, 2, -39, 9, 37, -1, -45, 38, -55, 63, 0, -48, 35, 8, -11, -5, -2, -62, 69, -11, -7, -4, 22, 9, -9, 32, 17, 23, -56, 11, 54, -75, 17, 15, -64, 56, -11, 27, -40, -43, 87, -41, -65, -12, 80, 12, -38, 76, -26, -80, 63, 76, -86, -24, 85, 35, -106, 14, 56, -51, 27, -23, 10, 20, -8, -32, -35, 3, -29, 14, 54, 39, -25, -15, 47, -59, 17, 29, -95, -6, 38, 59, 47, -24, -56, 41, 7, -52, 56, -47, -80, 62, 17, 43, -26, -80, 8, 25, 17, -38, 41, 66, 21, -75, -37, 68, -25, -15, -35, -7, 63, 4, -36, 19, -22, 19, 38, -13, -8, -38, 48, 21, -87, -20, 63, -25, -6, 54, 1, 6, 36, -46, -13, 54, -12, -51, 12, -37, 20, 69, -45, -2, -38, 51, -7, -59, 69, 27, -51, -52, 13, -24, 61, 15, -41, 14, 8, -29, -42, 10, 89, -28, -37, 98, -88, -27, 25, 15, 47, -66, -2, 2, 15, 74, -78, 28, 32, -120, 58, 69, -57, -60, 69, 1, -44, 27, 14, -34, -23, 85, -21, -44, 74, -36, -80, 100, 23, -57, 28, -41, 10, 1, -36, 28, 48, 19, -53, -27, 31, -17, 21, 86, -79, 5, -28, 9, 10, -31, 88, -14, -37, -25, -38, 14, 27, -7, 6, -60, 72, 9, -100, 85, -10, -2, -1, -48, 13, 35, 13, 25, 42, -56, 17, -18, -53, -6, -28, 46, 74, -53, -55, 37, 8, 0, 31, 36, 14, -74, 0, 82, -68, -76, 35, 35, 7, 12, -12, 44, -42, -88, 69, 85, -31, -20, -43, 26, 60, -72, -11, 22, -14, 21, 37, 17, -71, -21, 76, -81, 18, 53, 3, -47, -24, 37, -9, -15, 48, -2, -82, 4, 19, -8, -43, 99, 58, -85, 39, 3, -24, 1, 26, -15, -92, 90, -21, -49, 46, 31, 2, -47, -1, 1, 17, -48, 40, 6, -62, 90, -18, -30, 73, 0, -19, -61, 10, 36, -35, 27, 37, -35, -79, 65, 36, -58, 22, 13, 23, -42, -40, 23, 0, 49, 4, 17, 22, -45, -69, -18, 23, 3, 62, -15, -83, 42, 11, 20, 56, 0, -43, 4, -38, -12, 49, -24, 61, -40, -97, 85, 5, -46, 86, 26, -89, -1, 65, -65, -68, 90, 4, -45, 5, -43, 49, 10, -19, 61, 51, -56, -29, 29, -77, 47, -5, -25, 25, 34, 45, -73, 8, 48, 12, -20, -11, -55, -22, 32, -30, 24, -9, -23, 91, -27, -43, 28, -17, 69, -22, -55, 12, 37, 62, -62, -23, 58, 20, -1, 1, -25, -53, 7, 23, -39, -9, -9, -2, 60, 1, -9, -29, 11, -11, -73, 99, 31, -43, -6, -11, 44, 26, 0, -7, -1, -43, -35, 55, -22, -32, 36, 40, 25, -68, -21, -13, 10, 57, -18, -17, -30, -26, 42, 73, -61, -7, 59, -7, -31, -61, 3, -10, 56, 94, -18, -36, -39, -30, -3, 29, 23, 31, -18, -38, -36, 48, 37, -20, -5, 41, -41, -36, 13, -1, 37, -47, 14, -38, 57, 70, -97, -47, 56, 91, -68, -49, 54, -18, 10, 27, 34, -56, -29, 17, -7, 46, -47, -58, 23, 59, -39, -15, 23, -25, -14, 38, 40, -23, 23, 7, -66, 38, 46, -7, 17, -1, -38, -42, 3, -30, -11, 18, 3, 51, 11, 19, -12, -32, 69, 6, -62, -61, -7, 51, 2, -21, -21, 43, 63, 2, -60, 19, 38, -14, 32, -60, 8, -27, -11, 105, -80, 1, 8, -54, 47, 20, -34, 32, 9, -77, 41, 34, -47, 37, -27, -22, 12, -47, 23, 54, 65, -38, -15, 10, -31, -6, 63, -46, -30, 77, -79, 24, 52, -71, -3, -31, 60, 69, -109, -39, 105, 20, -3, -31, -31, -29, 32, 69, -77, -31, 32, -13, 40, -4, 0, 8, -11, 63, -41, -18, 5, 12, 2, -48, -56, 85, 30, -106, 44, 31, -35, 37, -35, -38, 95, 20, -69, 40, -23, -10, -12, -10, 87, 2, 7, -5, -81, 18, 34, -9, 0, -69, 5, 91, -29, -47, 66, -2, -19, -23, 31, 58, -9, 18, -72, -4, 37, -28, 13, 15, -41, -1, 26, -68, 26, 10, 15, 59, -82, -37, 48, 2, 4, -54, -15, 85, 6, -60, -4, -14, 25, 28, -70, 39, 23, -26, 9, 60, -32, -86, 77, 10, 27, -30, -32, 53, -20, 8, -24, 31, -54, 26, 38, -73, 82, 21, -74, -21, 71, 7, -34, -11, 34, 27, -90, -29, 0, 34, 10, -54, 60, 62, -20, -3, -57, -29, 26, 12, 66, 4, -65, 32, 28, -28, -15, 0, -8, 17, -19, -45, 27, 30, 53, -47, -27, -37, 9, 64, -22, 20, 30, -52, -9, 32, -76, 22, 92, -48, -53, 69, -46, -7, 80, -15, -14, -48, -14, 89, -53, -32, 43, -28, 21, -37, 38, 82, -75, -39, 32, 34, -20, -48, 6, -52, 75, 19, -26, 56, -8, -58, -10, 80, -69, -40, 64, 2, 23, -59, -17, 81, -5, 25, -35, -75, 6, 2, -11, 22, 54, 20, -31, -56, -27, 62, 4, -82, 85, 87, -28, -12, -64, -18, 44, -43, 54, -23, -14, 75, -87, -7, 22, 41, -6, -31, 80, -23, -6, -23, -90, 46, 87, -31, -29, 62, 30, -27, -2, 24, -31, -10, -11, 18, -52, 12, 89, 0, -102, -15, 75, -78, -44, 78, 76, -55, -42, 44, 55, -73, 1, 78, -29, 0, -44, -39, 57, -11, -65, 57, -10, 13, 23, -18, 35, -30, 14, 9, -28, 21, -4, -85, 59, 37, -7, 45, -109, -27, 68, 37, 9, -41, 26, 1, -45, -19, -35, -6, 58, -9, 27, 71, -86, -37, 48, 56, -66, -46, 66, 12, -21, -70, 64, 10, -34, 81, -78, -5, 27, -9, 53, -75, -24, 56, 14, 21, 14, 3, -77, -18, 14, -48, 30, 17, 24, -27, -32, 64, 35, -77, -7, 9, -37, 37, 0, 63, -14, -53, 54, 7, -36, -24, 43, 45, -81, -24, 65, 45, -44, -8, 26, -31, -55, 38, 97, -32, -80, -26, 34, 43, -12, 5, 55, -29, -47, -35, 34, 21, 21, -22, -55, -14, 41, 80, 8, -17, -39, -13, 25, 24, -22, -55, -5, 30, -19, -17, 1, -9, 45, 32, -54, -55, 38, 89, 3, -8, -37, -53, 35, -39, 14, 69, -53, -30, 56, -26, -47, -1, 49, 69, 22, -61, -78, 15, 59, -3, -21, 60, 6, -65, -15, 62, -35, 24, 40, -8, 11, 1, -38, -88, 78, 63, -19, -64, -56, 37, -2, -11, 12, 71, -38, -53, 9, -26, 54, 46, -7, -59, 19, -3, -14, -17, 39, 83, -109, -7, 72, 14, -28, 34, -48, -63, 100, 20, -17, -65, -51, 91, 7, -35, 52, -28, 22, 37, -32, -13, -3, -43, 37, -7, -43, 23, -29, 17, -24, -23, 95, 45, -95, -22, 80, -58, 27, 47, -13, 7, -21, -40, -11, -13, 34, 19, -41, 79, -56, -51, 42, 28, 20, -54, 43, -25, -28, 17, -31, 57, -6, -22, -8, 7, 45, 48, -27, -18, 3, -19, -9, -38, 29, 66, -49, -21, -28, 41, 31, -83, -5, 54, 55, 11, -86, -11, 97, -27, 4, -22, -62, -2, 44, 17, 6, 0, -24, 0, -18, -40, 72, 59, -79, 14, 12, 4, -32, -11, 48, -22, 14, 39, -58, -18, 49, -36, -28, 12, 73, -46, -8, 9, -46, 37, 24, -19, -74, 1, 70, -2, -38, 32, 56, 14, -65, -18, 14, 11, -30, -45, -7, 73, 85, -66, -31, 21, 6, 49, -76, -7, 3, 4, 91, -42, -45, 3, 48, -31, 7, 7, -13, -10, -71, 44, 92, -25, -86, 20, -12, -27, 64, -22, -40, 37, 23, 13, 58, -57, -25, -18, 25, 68, -15, 26, -65, -41, 30, -38, 40, 15, -28, 28, -18, 34, -40, -13, 6, -14, -11, -25, 70, 29, -47, 52, -45, -5, 85, -102, -37, 36, -10, -13, -2, -22, 100, 19, -59, 19, 0, -20, 35, -27, 8, 17, 6, -32, 4, 15, -71, 103, -11, -86, 21, 49, 52, -24, -41, 24, -14, 9, 42, -21, -5, 36, -22, 2, -37, -59, -1, 57, 11, 10, 51, -69, -59, 55, 8, -76, 52, 51, 26, -72, -13, 46, -21, 36, 20, -40, -52, 27, -34, -6, -15, 74, 7, -35, 76, -32, -72, -37, 24, 48, -23, -56, 94, 4, 1, -10, -51, 51, 41, -22, -21, 25, 21, -21, -47, 44, 23, 13, -62, 14, 5, -78, 89, 8, -89, 30, 91, -75, -4, 6, -24, 81, -53, -21, -3, -52, 58, 36, 1, -11, 31, -1, -97, 57, 64, -34, -10, 2, -22, 37, -4, -15, -18, -26, -5, 2, 5, -46, 42, 88, -40, -70, 57, 19, 0, 29, -9, -35, -22, -10, 62, -12, -11, -11, -66, 56, 39, 32, -53, -70, 72, 29, 24, -57, -85, 18, 32, 8, -27, -10, -14, 42, 9, 19, 82, -83, -38, 74, -31, 48, -49, -55, 37, 27, 20, -29, -4, -28, 2, 29, 12, -38, -27, 38, -4, -20, 34, 29, -9, 7, 18, -6, -43, -62, 35, 15, -32, -23, 70, 70, -111, 45, 9, -73, 76, 6, 34, -65, 0, 36, -36, 14, -23, 52, 29, -7, -61, -23, 20, 37, -15, -71, 32, 30, -42, 48, 51, -78, 46, 8, -10, 65, -58, -90, 15, -6, 29, 27, -69, 32, 40, 5, 46, -71, -31, 75, 8, 19, -61, -57, 56, 8, -12, -43, 40, 78, -110, 2, 18, -66, 12, 9, -19, 45, 11, -24, 39, 43, 1, -9, -15, -46, 19, 3, -6, -12, -32, 26, -13, -2, 60, 18, 32, -64, -3, 74, -12, 18, -35, -102, 63, 64, -90, -43, -2, 34, 20, 38, -12, -65, 28, 55, -1, -62, -48, 104, 11, -78, 20, -5, 51, -30, -73, 80, 11, -78, 42, 23, -58, -14, 34, -12, 30, 56, -78, 31, 86, -38, -17, -41, 29, -14, 17, 28, -78, -7, -2, 49, 3, -4, 70, -60, -13, -6, 20, -1, -85, 66, -3, -26, 29, 29, -19, -27, -26, 32, 0, -48, -1, 72, 0, 5, 78, -74, -54, 0, 6, 35, 28, 31, -62, 8, -26, 13, 92, -29, 34, -82, -51, 29, -19, 71, 38, -14, -72, 32, 13, -70, -14, 11, 1, -14, 19, 59, 21, -36, -52, 52, -3, -24, 85, -64, -15, 55, -30, -37, 52, -21, -6, -19, -13, 106, -61, -61, 89, -24, -24, -27, 17, 49, -35, 21, 30, 4, -11, -34, -34, 46, -4, -38, 47, -57, 31, 6, 1, 1, -29, 53, -22, -37, 31, -9, -63, 82, 15, 27, -53, 11, -2, -35, 62, -40, 8, -19, -12, -24, 37, 44, 0, 55, -85, -41, -2, 35, 56, -1, -53, -62, 52, 11, 13, -47, 3, 59, 35, -68, -26, 115, -80, -24, 79, -23, -40, -45, 71, 35, -72, 18, -11, -47, 51, -5, 1, 48, -60, -30, 46, -23, -3, 79, -9, 7, 52, -97, -20, 83, -56, -43, 63, -4, -68, 13, 86, -23, -28, 47, 30, -80, -46, 21, -36, 94, -7, -9, 29, -44, -42, 53, 42, -48, 43, -57, -17, 71, -42, -34, 21, 10, 34, -45, 8, 73, -34, 7, -42, -43, 55, -29, -30, 99, -31, -44, 81, -17, -34, -24, 49, 32, -82, 6, -13, 48, 39, -29, 7, 17, -45, -80, 29, 74, -11, -69, 36, 62, 26, -3, -68, -31, 75, 10, -43, -45, -10, 14, 26, 45, -9, -8, -35, 39, -26, -46, 89, 9, -55, -13, 26, -10, -4, 60, -48, 2, -10, -12, 89, -98, 6, -3, -13, 58, 8, -56, -7, 110, -43, -66, 42, 54, 35, -105, 6, 5, -40, 77, -7, 38, -52, -66, 24, 54, -28, -21, 57, -42, -9, 9, -5, -27, 9, -22, 31, 19, -82, 48, -3, -11, 70, 39, -46, -9, 70, -62, -6, 51, -99, 10, 66, -61, 56, -19, -94, 25, 48, 53, -17, -47, -48, 89, 13, -61, 91, -68, -18, 7, -40, 90, -6, -57, 13, 78, -71, -25, 17, 35, 2, -80, 47, 46, -4, -30, 27, 9, -5, -11, -26, -22, 26, 36, -46, -48, -2, 21, -23, 69, 8, -39, 45, 0, 32, -52, -27, 75, 8, -9, -1, 30, -69, -63, 78, 11, 15, -3, -66, 32, -39, -3, 100, -10, -52, -60, 51, 34, -59, 51, -10, -27, 9, 31, -4, -68, -19, 79, -15, -8, 69, -17, 22, -3, -57, -12, 29, -39, -36, 54, 81, -74, -35, 69, 25, 0, 9, -13, -58, -26, 14, 23, 34, 23, -32, -58, -46, 57, -3, -58, 47, 63, -53, -41, 62, -23, 60, -41, -39, 20, 12, 43, -57, 1, 0, -11, 0, -10, 66, 30, -37, -6, -37, 21, -4, 19, 51, -48, -32, 48, 1, 15, 0, -31, -4, -52, -29, 31, 0, 22, 27, 37, -45, -6, 34, -46, -13, 8, 76, -60, -46, 39, 20, 27, -75, 41, 44, -22, -5, 9, 47, -121, 49, 23, -36, 25, -48, 48, 30, -26, -19, -28, 6, 44, -57, 44, -2, -72, 55, 54, -20, 4, 2, -89, 31, 38, -47, -32, 13, 56, -42, 39, 71, -106, -24, 34, 4, 40, -28, -52, 14, 40, 6, 25, -25, -28, 70, -51, 32, 9, -88, 36, -6, 6, 35, 25, -64, -11, 104, -49, -69, 82, -10, 1, -24, -37, 36, -19, 7, -13, 38, 19, -62, -42, 44, -1, 43, -21, -28, 78, -35, 18, -22, -15, 23, 11, 9, -43, 23, -19, 17, 63, -48, -81, 65, 12, -3, -32, 19, 1, -46, 60, -1, 1, 17, -70, 22, 59, -92, 17, -1, 9, 12, -21, -8, 36, -8, 2, -6, 11, -17, 9, 77, -69, -46, 8, 58, 37, -23, -34, 59, -51, -85, 60, 39, 22, -8, -24, -30, 11, 80, -32, -66, -15, 57, 11, 17, -40, -74, 9, 59, 19, -90, 25, 64, -49, 32, 32, -102, 11, 89, 45, -39, -83, 17, -3, 48, -12, -23, 18, -1, 56, -14, -69, 39, 43, -56, 59, -22, 2, -43, -49, 22, -44, 69, 61, -68, -8, 92, -37, -113, 94, 7, -40, -9, 4, 70, 14, 14, -46, -59, 35, -11, 14, 77, -85, -30, 41, -49, 61, 21, -92, 13, 18, -1, -27, -29, 40, 76, -69, 4, 74, 0, 36, -80, 9, 61, -124, 47, 49, -58, -8, -48, 68, -17, 7, 94, -51, -38, -44, 10, 71, -45, 28, -21, -46, 111, -54, -95, 74, -12, 20, 13, 11, 55, -69, 45, -20, -55, 69, 30, -89, -75, 96, 64, -92, 18, 45, -8, -45, 2, 4, 0, 92, -103, 4, 44, -14, 63, -51, -52, 72, -31, -36, 82, 18, -80, 17, -1, -27, 89, -102, -2, 100, -5, -24, -85, 34, -2, 0, 77, 0, -85, -10, 90, -79, -5, 22, -68, 34, 60, -3, -26, 49, -21, -55, 71, 5, -38, -42, 3, 26, -32, 1, 17, -37, 63, 23, -1, -28, -68, 75, 58, -40, -44, 37, 14, -73, 40, 57, -40, 11, -40, -45, 41, 28, 8, 0, -52, -29, 46, 42, -22, 15, 43, -8, 0, 14, -76, -1, 74, -30, -36, 44, -52, -82, 60, 51, -42, -5, -3, 48, -19, -39, 1, 21, -10, 9, 24, -87, 95, 46, -21, -18, -27, 40, -30, -23, 35, 4, -24, 0, -26, 48, 22, -76, -30, 62, 87, -78, -34, -4, -29, 34, 44, -25, -52, 32, 97, -51, -29, 78, 14, -30, -53, 11, -17, 29, -34, 19, 34, -59, 19, 9, -7, 19, 45, -42, -6, 19, 13, -64, -5, 97, -31, -48, -40, 25, 96, -76, -3, 85, -113, 37, 28, -54, 27, 15, -25, -6, 37, 7, -44, -54, 17, 55, -36, -45, 14, 45, 64, 7, 2, -32, 13, -9, -83, -25, 17, -9, 11, -5, 54, 32, -79, -26, 89, 35, -9, -22, -62, 25, 75, -18, -29, 5, -74, 45, 46, -57, 2, 20, -29, 1, -10, -35, 86, -3, -82, 107, -14, -47, -9, 37, 93, -93, -75, 72, 51, 24, -61, -100, 73, -11, -4, 23, -24, 34, 46, 22, -3, -42, -47, -32, 48, 30, -65, 25, 26, -15, -1, 12, 45, -13, -37, 27, 4, -3, -11, -31, 20, 11, -17, -37, 1, 90, -39, 0, 30, -83, 43, 4, -35, 87, -26, -73, 5, 17, 41, 10, 25, -53, -66, 70, 21, 7, -14, -60, 5, 60, -2, 29, -39, 2, -10, -36, 91, -53, -11, -12, -1, 6, -6, -10, -41, 78, 2, -31, -13, 64, -2, -103, 14, 20, 58, 36, -58, -70, 86, 35, -8, -4, -27, -25, -25, 48, 53, -69, 19, 38, -81, 22, 23, 25, -15, 7, -9, 8, -25, -25, 75, -51, -12, 64, -7, -44, -10, 42, -3, -36, -10, -9, 48, 48, -35, -66, 9, 14, -23, 9, 34, 5, 27, -30, -58, 11, 64, 43, -90, -48, 18, 74, -10, 7, 27, 0, -14, -94, 44, 68, -40, 35, -31, -81, 86, 18, -31, -37, 35, 54, -28, -22, -27, 0, 35, 2, 12, 13, -64, 31, 52, -45, 17, -52, -18, 46, -71, 56, 40, -22, 12, 22, 8, -21, -35, -18, -1, 19, 56, -79, -12, 27, -11, 48, 25, -64, -37, 38, 37, 7, -40, 0, -15, -45, 40, 57, -21, -5, 0, 39, -9, -99, 88, -25, -8, 29, -40, -9, 47, 15, -87, 38, 19, 35, -25, -65, 82, 24, -25, 31, -59, -45, 7, 17, 0, 49, -37, 1, 42, -36, 43, 7, 0, -6, 6, 10, -91, -32, 113, -63, -14, 24, -24, 5, 37, 62, -61, 29, -4, -63, 38, 23, 2, -63, -44, 1, 75, 6, 5, 5, -10, 69, -98, 9, 59, -90, 0, 59, -8, -20, 20, -27, 4, -4, -22, 63, -56, -58, 70, 26, -9, -2, -37, -9, 23, 7, -3, -12, 36, 0, -9, 51, -69, 27, 37, -30, 71, -75, -58, 60, 15, -61, 37, 19, -65, 15, 59, -9, -41, 17, 38, -52, -7, 115, -63, -71, 10, 40, 26, -87, 65, 12, -39, 20, -71, 0, 100, -22, -73, 43, 17, 55, -21, -32, -36, 22, 72, 22, -77, -59, 39, 48, 0, -74, 52, 44, -37, -45, -21, 97, -24, -64, 0, 47, 43, -69, -40, 29, 22, -22, 49, 61, -61, -61, 26, 11, -37, -11, 35, -23, 22, 55, 26, 19, -1, -12, -21, -42, 48, -42, -53, 24, -18, 40, 52, 23, -9, -79, -34, 9, 5, 17, -60, 59, 44, -30, -39, 6, 71, -28, 3, 1, -65, 48, 18, -65, 38, -26, 6, 63, -66, -45, 68, 26, -8, 29, -37, -15, 38, 15, -3, -63, 35, 45, -7, -8, -95, 65, 85, -25, -52, 0, -28, -3, 29, -29, 42, 44, -34, -42, -1, 8, 23, -70, 59, 14, -37, 20, -5, 24, -74, -7, 49, 48, 38, -45, -53, -37, 19, 12, 29, 57, -8, 23, -40, -71, 12, 3, -44, 71, 49, -47, -6, -39, 18, 27, -23, -20, 47, -25, -19, 87, -36, -58, 45, 0, 6, -28, -35, 26, -18, 17, -29, -4, 19, 22, 17, 11, 24, -8, -7, -14, -34, -38, 35, 76, -32, 35, -35, -73, 4, 57, -9, -28, 2, 13, 85, -14, 10, -64, 30, -7, -70, 115, -36, -24, 23, 0, 6, -63, 14, -24, 11, 71, -61, -38, 32, 38, -25, -22, 77, -19, -74, 68, 58, -75, -6, 53, -68, -21, 103, -60, -31, 59, -79, 68, 9, -55, 71, -8, 18, -49, -9, 30, 0, 38, -10, -54, -32, 73, 32, -66, -38, -20, 0, 0, -2, 85, 31, -48, -27, 24, 0, 52, -49, -56, 119, -43, -85, 51, 85, -91, 2, 76, -62, 22, 2, -47, -56, 83, 1, -19, 19, -58, 74, -6, -35, -20, -10, -3, 18, 52, 22, -70, -8, 81, -12, -21, 37, 32, -82, 10, 74, -81, -21, 9, 54, -39, -57, 113, 19, -32, 1, -54, -70, 54, 31, -12, 11, 20, 5, -60, -18, 26, -43, 88, -24, -31, 63, 12, 1, -22, 47, -37, -80, 0, 89, -47, -40, 53, -48, 4, -4, 44, 40, -73, -10, 72, 24, 0, 4, -62, -40, -34, 57, 8, 28, 53, -113, 3, 62, -2, -19, 1, -36, -9, 92, 28, -35, -37, -30, 26, 55, -34, -14, -17, 1, 85, -56, -61, 82, 36, -8, -91, 25, 44, -83, 79, -40, -58, 58, 23, -61, 38, 26, -99, 49, 3, -45, -7, 59, 13, 21, 0, 1, 3, -18, 26, -27, -53, -32, 36, 75, 45, -54, 13, -24, -2, 69, -65, -39, 14, -40, 11, 32, -35, 27, 62, -32, 1, -37, -61, 14, 70, 49, -95, -11, 30, 21, 53, -43, 9, -1, -57, 53, 54, -42, -85, 76, 0, -36, 17, -4, 34, 27, -59, -90, 55, 88, -6, -74, 52, 38, -60, 35, -25, -21, 0, 6, 21, -61, -13, 8, 25, 40, -45, -29, 109, -22, -63, -1, 54, 42, -6, -1, -20, -69, 19, 12, 22, 11, -60, 75, 46, -102, 1, 20, -10, -21, 29, 10, -86, 20, -1, 54, 36, -26, -64, 31, 62, -41, 32, 25, -92, 47, 2, -21, 91, -89, -95, 112, 8, -43, 77, -55, -9, 52, -31, -20, 28, 1, -31, 56, -1, -10, 20, -56, -40, 64, -22, -89, 45, -11, 28, 43, 36, -57, -66, 126, -60, -47, 105, -27, -71, 45, 51, -85, -11, 21, 8, -4, 21, -1, -60, 43, -36, 51, 78, -75, 5, 54, -29, -86, 65, -2, -42, 104, -61, -85, 95, -9, -19, 65, -17, -70, 0, 35, -42, -29, 34, 77, -34, -54, 75, 14, -12, -52, -21, 63, -18, -12, -12, 63, 9, -58, -28, -7, 20, -1, 21, -18, 10, 19, -64, -2, 40, 25, 10, -1, 18, -47, -14, -18, 10, 37, 0, 0, -13, -20, 39, 80, -35, -64, 53, -27, -10, 3, -32, 9, 0, -10, -8, 12, -11, 41, -13, 48, -22, -92, 47, 82, -26, -99, 68, 93, -64, -19, -19, 29, 70, -91, 20, 31, -42, 53, 4, -30, -57, -27, 69, 34, -36, -48, 45, 59, -9, -58, 18, -32, -39, 45, 29, 45, -56, 9, 25, 9, -10, -106, 64, 35, -83, 61, 68, -104, 2, 72, -25, -55, -65, 45, 69, -11, -3, 26, -43, -17, 80, -45, -46, 42, -3, 3, -24, -36, 10, 2, -46, 90, 8, -92, 13, 34, 81, -52, -42, 81, 20, -65, 4, 65, -22, -13, -38, -5, -10, 8, 92, -63, -10, 41, -21, -12, 23, 64, -52, -52, -46, 35, 14, -57, 57, 4, 1, 24, -26, -21, -5, -6, 21, 0, -51, 1, 75, 2, -25, 62, 30, -23, -91, 40, -7, 0, 28, -94, 66, 66, -56, 21, -9, -18, -36, 24, 99, -35, -37, -41, 55, 45, -47, -32, 45, 10, -30, 10, 31, -36, -39, 88, -86, -17, 106, -94, 5, 0, -49, 48, 43, 26, -41, -54, 5, 30, -28, -4, -1, 20, 64, -58, -20, 14, 21, 3, 25, 10, -98, 61, 61, -23, 15, -2, -20, 9, -72, -38, 98, -7, -99, 52, 19, -52, 90, 3, 1, -31, -91, 0, 78, 63, -58, -30, -10, -40, 83, -6, -29, 8, -55, 29, 94, -39, -81, 77, 56, -41, -70, 43, 58, -56, -35, 77, 22, -58, -7, 24, 0, -11, 25, -10, -38, -32, 46, 41, -72, 22, 36, 6, 6, 4, -52, -11, 73, -23, -42, 20, 42, -2, -43, -7, 48, 29, -42, -15, -6, -53, -12, 81, 47, -98, -15, 9, -21, 8, 32, 15, 28, -19, -65, 35, 71, -5, -87, 58, -32, -19, 56, 13, -22, 10, 27, -88, 68, -40, 8, 38, -93, 21, -13, 68, 8, -27, -30, -11, 91, -1, -82, 7, 87, -37, -66, 48, 66, -44, -25, 57, -42, -81, 70, 43, -66, -37, 92, -22, -74, 104, -10, -31, -9, 0, 34, 0, -28, 0, 8, -49, 0, 13, 72, -45, 1, 1, 3, 66, -43, 3, -9, 23, 29, -49, -18, -39, 25, 52, -63, -25, 20, 40, 28, 11, -47, -28, 7, 36, -48, -1, 99, -49, -75, 57, 40, -100, 59, 44, -35, 37, -66, -21, 62, -59, 41, 20, -95, 70, 46, -24, -69, -18, 14, 48, 80, -32, -69, 1, 1, -7, 1, -31, 56, 12, 26, -14, -65, 85, 28, -75, -12, 72, 12, -62, -73, 56, 44, -57, 14, -19, 29, 35, -36, -45, -5, 46, 10, 15, 23, 35, -82, -64, 2, 62, 61, -83, -43, 19, -20, 75, 31, -32, 58, -45, -76, -14, -9, 59, 19, -14, 63, -41, -71, 25, 1, 15, 49, 35, -58, -15, 70, -53, 10, 74, -81, -18, -9, -35, 90, -29, -48, 30, -41, -11, 76, -26, -46, 70, 30, -6, -36, -15, 62, -21, 9, -24, -92, 59, 95, -40, -65, 54, 39, -57, 17, -40, 13, 97, -76, 15, -45, 9, 22, -87, 1, 76, -1, -45, 32, 54, -56, -2, 37, 4, 3, -89, 92, -2, -25, 75, -25, -70, 18, 12, -14, 13, -25, 23, -25, 35, 14, -70, 46, 13, -44, 47, -20, -22, 0, 13, 28, -54, 10, 65, -49, 11, 0, -73, 30, -25, -15, 97, -5, 0, 22, -111, 13, 85, 1, -9, 29, -76, -56, 55, 27, 12, -29, 32, -12, -29, 46, 11, -60, -52, 76, 1, -60, 56, 42, -52, 31, 44, -46, -63, 46, 62, -63, -45, 34, 69, -56, -66, 107, -25, -8, 23, 6, -20, -55, -6, 63, -28, -13, 116, -85, -23, 1, -11, 11, 23, 68, -72, -17, 20, -25, 29, -49, 24, 72, -13, 4, -76, -58, 87, 8, -68, 1, 19, 2, 36, 13, -44, 28, 19, -44, -31, -26, 51, 45, -14, -13, 0, 46, -57, 23, 21, -28, -4, -64, 45, 69, 28, -29, -76, 3, 90, -56, 8, -3, -29, 45, -13, 58, -42, -81, 15, 14, -17, 47, 60, -12, -57, -28, 30, -2, -29, 56, -27, -55, 103, 13, -76, 40, -15, -42, 46, -61, 38, 30, -62, 11, 49, 57, -41, -80, -24, 63, 23, -41, 21, -4, -55, 53, 55, -19, -60, 47, 32, -91, 15, 0, 35, 54, -93, 41, 11, -66, 94, 25, -14, -59, -54, 57, -23, -6, 66, -46, -53, 91, 22, -30, -25, -9, 18, 29, -29, -43, 82, -22, 0, -35, 2, 35, -7, 46, -57, 25, -1, -75, 54, 71, -43, 1, 17, -47, 18, -51, 17, 75, -71, -47, 42, -7, 32, 63, -91, 25, 17, -5, 2, 14, -20, -106, 55, 58, 28, -2, -2, -64, -58, 52, -14, 11, 30, 3, -34, 27, 65, -15, -9, 13, -43, -81, 7, 79, 72, -81, 14, -2, -70, 18, -4, 0, 0, 51, -28, -60, 47, 58, -35, -5, -2, -28, 4, 6, 88, -31, -55, 60, -27, -64, 53, 19, -55, 62, 9, -76, 3, 2, 12, 27, 1, 8, 24, 24, -54, 18, -38, -4, 76, -74, -10, 53, 8, -7, -28, 5, -44, 29, 44, -74, -10, -34, 61, 21, 6, 72, -32, -77, -37, 92, 36, -37, 12, -30, 6, -41, -31, 60, 43, 24, 9, -59, -13, 38, -71, -40, 24, -23, 80, 47, -71, -41, 11, 100, -21, -66, 59, 53, -32, -88, 57, -1, -12, 47, -29, -4, 3, -40, -58, 70, -14, -66, 102, 58, -25, -79, 17, 108, -105, 12, 41, -44, -30, -54, 57, 32, -9, 6, 0, -47, 30, 35, -49, 40, -31, -55, 14, 63, -6, -39, 24, -24, 25, -9, 59, -4, -91, 104, -32, -60, 95, -10, 8, 38, -43, -24, -19, -51, 70, 70, -98, 13, -9, -14, 31, -60, 45, 23, 5, 37, 4, -85, 36, 26, -94, 97, -1, -48, 64, -11, -90, 44, 0, -80, 62, 48, -12, 20, 20, -32, -25, 58, -43, -32, 44, -36, 42, -45, 11, 44, -8, 17, -38, 27, 18, 1, 11, -72, -25, 54, 5, -1, -32, 6, 26, 27, -32, -76, 47, 75, 1, -88, 22, 66, -10, -43, -55, 28, 20, -65, 77, 9, -52, 61, -75, -8, 38, 29, 8, 12, -4, -77, 11, 48, 42, -73, -10, 8, -42, 37, -47, 75, 37, -24, 53, -66, -45, -25, 54, 64, -90, 22, 73, -7, -53, 22, -19, -13, 53, -13, 23, -88, 45, 8, -36, 88, -65, -44, 74, 7, -31, 48, -8, -88, 46, 17, -38, -19, -5, 17, 18, 40, -74, 4, 29, -17, 5, 9, -8, -52, -1, 102, -27, -65, -2, 70, 0, -64, 25, 49, 54, -7, 9, -45, -72, 34, 64, -22, 14, -53, 17, 31, -15, -34, -75, 15, 38, 21, 6, 30, -31, 26, 15, -37, -39, 12, 32, -62, 62, 57, -103, 24, 70, -92, -42, 87, 53, -92, -20, 68, -38, -3, -8, -51, 51, 6, -55, 90, 26, -25, 8, 14, 21, -88, -21, 71, 19, -9, 30, -11, -43, -48, 10, 5, -51, 60, 74, 2, -11, -36, -41, 62, 46, -52, -75, -13, 64, -20, -32, -17, 64, 60, 1, -24, -7, 0, -66, 34, -11, -31, 3, 34, 7, -4, 43, -24, -37, 26, 0, -73, 79, 70, -121, 39, 14, -85, 4, 62, 7, -55, 70, -39, 28, 65, -65, 26, 43, 1, -55, -57, -30, 38, 68, -23, -54, 0, 64, -3, 27, -46, -54, 107, 0, -37, 10, 17, -14, 14, -31, 12, -15, -100, 111, -10, -30, 43, 11, 34, -66, -39, 65, -9, 1, 23, -10, -55, 22, 53, -59, 49, 4, -91, 45, 2, -18, 35, 20, -9, -64, 11, -19, 9, 25, -43, 22, -6, 0, 36, 4, 44, -6, -17, -55, 14, -17, 26, 51, 5, -9, -98, 55, 82, -78, -7, -25, 37, 1, -3, 26, -62, 12, -12, 61, 11, -34, -29, 27, -35, 5, 31, 10, 0, 12, -45, 18, -2, -22, 90, -109, -27, 78, 56, -58, -85, 48, 5, 40, 49, -87, -20, -11, 12, 54, 49, -62, -66, 19, 53, -13, 26, -2, -96, 48, -13, -26, 43, -13, -44, 111, -13, -74, 81, 42, -22, -4, -20, 2, 57, -83, -59, 14, -4, 41, 73, -64, 0, 2, -44, 54, -10, -17, 27, 8, 7, 12, 5, -60, -5, 93, -83, 4, 14, -1, 48, -8, 14, -87, 18, 52, -80, 48, 44, -61, 2, 2, 5, -19, -13, 73, 8, -2, -34, -52, 5, 60, 71, -102, -86, 66, 78, -60, -36, -12, 48, 98, -23, -24, -81, 17, 2, -45, 46, 25, 7, 23, 49, -77, -88, 59, -27, 35, 34, -60, -17, 38, 24, -80, 51, 25, -9, 18, -32, 63, 0, -73, 73, -24, 13, -31, -5, 15, -76, 44, 18, 63, -47, -17, -14, -22, 18, -42, 13, 29, 10, -3, -42, 37, 27, -14, 61, 38, -87, -61, 100, 0, -20, 39, 0, -9, 8, -6, 4, -44, -76, 47, -5, -8, 8, -40, 83, 1, -58, -12, 29, 64, -40, 13, -14, 6, 19, -65, 48, 17, -14, 39, -71, -15, 74, -71, -22, 61, 37, -36, -3, 71, 6, -98, -25, 12, -28, 38, -4, 25, 20, -62, -21, 93, 38, -37, 10, -34, -79, 35, 73, 20, -59, 24, 4, -6, 62, -19, -32, 6, -38, -39, 82, -53, -24, 36, -60, 61, 48, -43, -1, -40, 4, 85, -61, -44, 48, 39, 8, -28, -12, -7, -12, 38, -4, -9, 55, -54, -8, 20, -66, 45, 73, -6, 13, -42, -62, -25, -3, 78, 23, -28, 58, -63, -31, -4, 3, -5, 37, 12, -35, 22, 0, -24, -47, 0, 54, 95, -57, -39, 2, 6, 2, -36, 23, -5, 13, 53, -53, 32, 15, -9, 25, -40, -49, -27, 47, 41, -30, -24, 55, 42, -3, -53, 19, 57, -57, -11, 39, 14, -54, -68, 23, 38, -9, 25, 53, -90, -12, 20, -57, 3, -9, 60, 56, -82, 57, -9, -19, 24, -39, 57, -45, -19, 1, -24, 17, 56, -38, -54, 73, -4, -5, -32, 34, 91, -9, 0, -87, -23, 108, -56, -18, -12, 25, 36, -95, 83, 22, -91, -4, -14, 55, 38, -29, -51, 12, 97, -20, -3, -46, -35, -8, 32, 42, -86, 36, 30, 2, 39, 6, 20, -106, -10, 94, 32, -86, -87, 115, 22, -64, -23, 34, -10, 13, 2, -64, 53, -35, 51, 25, -81, 17, -5, 63, 36, -69, 8, -23, -48, 45, -12, -46, 31, 64, 52, -46, -2, -17, -43, 24, 6, 24, 37, 18, -53, -51, -44, 88, 23, -104, 3, 54, 2, -3, 31, -75, 61, 15, -97, 17, 40, 2, -52, 73, 89, -94, -64, 87, -23, 7, -23, 4, 52, -98, 27, 89, -61, -14, 68, -37, -6, 45, 40, -97, -46, 70, -61, -5, 64, -44, 10, -3, -42, 68, 70, -65, -4, 4, 17, -6, -99, -2, 89, 41, -102, 29, 18, -29, -9, 66, 47, -20, 23, -26, 14, -22, -89, 68, 57, -23, -63, -41, 82, 2, -82, 42, 44, 23, -62, -46, 127, -76, -44, 107, -36, -13, 0, -14, 66, -9, -40, 22, -10, -20, -1, -13, 47, 19, -59, 19, -5, -12, -21, -56, 106, -15, -12, 63, -109, 55, 17, -112, 93, 58, -2, -34, -46, 18, -48, 0, 97, 23, -91, 0, 3, -5, 96, -61, -72, 38, 46, 12, 6, 26, -22, 18, -82, -11, 56, -76, 22, 51, -53, 0, 24, -57, 56, 70, -61, 29, -21, -54, 52, -22, 34, 56, -114, 18, 103, -76, -51, 38, 68, -48, -47, 71, -55, -15, 39, -19, 20, 60, -78, -10, 61, -78, 65, 4, -97, 25, 10, -26, 64, 41, -27, 9, -17, -11, 29, -43, 24, 63, -5, 4, -76, -30, 51, -18, -65, 69, 74, -45, 17, 15, -38, -34, -36, 5, 61, -42, 11, 71, -51, -13, 20, -56, -26, 96, 22, 1, -39, -43, 88, -48, -37, -11, 35, -4, -53, 102, -48, -64, 52, 76, -48, -93, 45, 3, 4, 82, -15, -72, 42, 43, 22, -73, 11, 17, -92, 57, -5, -18, 15, -49, 46, 68, -60, -28, 60, 21, -59, 11, 64, -5, -20, 12, 32, -91, -69, 37, 80, 5, -36, 31, -40, -12, 70, -51, 5, -20, 7, 0, -40, 23, -49, 9, 69, 0, -17, 20, 18, 54, -81, -2, 45, 5, 10, -29, -82, 29, 97, -1, -54, -25, 25, 14, -38, -13, -12, -54, 56, 82, -51, -92, 108, 5, -83, 70, 4, 27, -23, -62, 79, 4, -64, 12, 32, -54, -37, 40, 88, -49, -47, 31, 30, -21, -62, -6, 52, 15, -60, 21, -10, -4, 39, -34, 4, 65, 31, -79, 4, 5, -28, 65, -11, 38, -36, -65, -14, 13, 89, -61, -11, 36, -28, 22, -7, 19, 17, -64, 36, 68, -65, 47, -51, -1, 10, -47, 65, 18, 8, -65, 51, -22, -3, 58, -94, -36, 82, -20, -21, 59, -58, -31, 71, 22, -10, -24, -44, 1, 23, -28, 46, 92, -95, -91, 89, 2, -25, 41, -65, -15, 88, -38, -38, 86, 0, -20, 47, -29, -18, 26, 27, -76, -5, 99, -55, 5, -57, 14, 94, -35, -103, 49, 57, -111, 73, 12, -82, 46, 32, -35, 29, 8, -55, 11, -19, -30, -7, 7, 30, 63, 36, -53, 7, 48, -65, -21, 27, -12, -5, 13, -46, 1, 44, -11, 27, -17, 22, -34, -81, 54, 41, -71, 42, 98, -58, -85, 66, 44, -79, 7, 19, -45, 63, 28, -106, 0, 95, 11, -12, 2, -88, 73, -18, -38, 59, 5, -30, -49, 87, -25, 5, 14, -77, 73, -19, -24, 97, -64, -66, 14, 34, 42, -30, 12, -44, -6, 9, -57, 9, 86, 32, -75, 47, 32, -95, -1, 41, -39, 61, -6, -41, 69, -14, 17, 3, -12, 13, -13, -51, -75, 93, 72, -35, -23, -27, 55, -53, -39, 109, -45, -42, 28, 10, 4, -69, 29, 88, -26, -95, 37, 76, -25, -7, -28, 11, -5, -38, 3, 72, 1, -73, 74, -18, -83, 25, 66, -52, -24, 28, 35, 40, -14, -25, -36, -12, 12, -2, -55, 102, -11, -17, 66, -17, -4, -74, -5, 79, -21, 2, 37, 0, -51, 0, -18, -22, 6, 27, 37, -21, -32, -15, 20, 40, 47, -14, -60, -49, 91, -8, -58, -9, -5, 7, -48, 81, 23, -51, 47, 21, -28, -24, 20, 31, -45, 4, 6, -40, 32, 45, -60, 0, 29, -41, 61, -32, -54, 86, 27, -74, -8, -30, 4, 77, -44, -19, 45, -24, 61, -19, -89, 30, 40, 46, -72, 20, 49, -66, 3, -29, -19, 32, 58, 10, -94, 6, 86, -37, -14, 3, 0, 64, -28, -82, 29, 34, 9, -56, 36, 69, -80, -29, -35, 76, 105, -107, 9, 40, -39, -8, -9, 53, 22, -38, -49, 58, -32, -74, 23, 43, 17, 24, -5, 8, -39, -87, 47, 57, -31, -25, 14, 0, 32, -20, -9, 24, 4, -2, -45, -31, 74, 55, -89, 9, 12, -27, 49, -38, 11, 47, 25, -61, -19, 42, -74, 32, 45, -24, -20, 13, 60, -8, -73, -18, 82, 5, 5, -1, -89, -39, 55, 77, -5, -9, -25, 27, -18, -87, -9, 81, 51, 14, -70, -57, 56, -32, -44, 81, 54, -66, 7, 2, 37, 22, -15, 28, -65, 11, 6, -61, 60, 61, -73, -34, 49, 12, -26, 9, 38, -38, 3, 0, -22, 21, 32, 9, 9, -103, 2, 62, -56, -11, 63, 1, -104, 74, 7, -57, 66, -7, 12, 13, -34, -39, -21, -4, 63, 64, -107, 13, 23, 7, -8, 1, 52, -90, 36, 38, -76, 18, 78, 0, -105, 34, 109, -98, 0, 4, -19, 39, -4, 18, -58, -38, 68, 11, -42, 44, -38, -15, 35, -11, -8, 25, -6, 18, 69, -85, -28, -10, 43, 27, -11, -37, -48, 96, -24, -49, -30, 70, 77, -34, 0, -73, -49, 46, 26, 20, -43, 14, 1, -8, 3, -7, 17, -7, 37, -48, 42, -18, -57, 88, 9, -69, 48, -18, -82, 25, 18, -3, -12, -11, 74, 72, -86, -62, 4, 55, 44, -36, -39, 45, 64, -38, -52, -7, -43, 74, 32, -22, 56, -2, -24, -25, -49, 1, 47, -42, 7, 70, -44, -7, 77, -61, -26, -8, -34, 71, 23, 29, -56, -106, 97, -15, -29, 25, -47, 62, -36, 10, 38, 17, 32, -100, -6, 75, -6, 18, 56, -92, -4, 31, -99, 49, 62, -31, 19, 47, -52, -45, 78, -22, -37, 41, -15, -65, 45, 51, -28, 30, -27, -80, 45, 93, -68, -72, 54, 58, -56, -2, -8, -60, 7, -15, 81, 46, -26, 9, 3, -58, -35, 58, 28, -72, -7, 13, -26, 15, 44, 78, -68, -71, 17, -23, 1, 43, -4, 57, -9, -37, 55, -42, 13, 39, -36, 4, -4, -43, 13, -22, -10, 69, 39, -92, 20, 27, -79, -4, 20, 104, -63, -23, 30, -65, 66, 5, 0, -25, -46, 97, 44, -105, -29, 61, 19, 44, -44, -72, 0, 58, -4, -11, 42, -79, 28, 39, -70, 64, 9, -25, 54, -31, -28, -49, 39, 13, -42, 40, -36, 45, 26, -102, 53, 83, -39, -13, 14, 24, 23, -96, -4, 15, 4, 14, -60, 36, 28, 2, -11, -48, -2, 18, 10, 60, -30, -36, -38, 36, 93, -74, -3, 5, -45, 47, -44, 53, 9, -29, 100, -103, 10, 72, -85, 18, 62, -10, -60, 4, -8, 17, 46, -11, -52, -30, 45, 4, 21, 6, -42, 0, 66, -72, 6, 21, -26, -10, -60, 95, 69, -72, -96, 78, 88, -69, -14, 60, -61, -74, 46, 17, 54, -18, -81, 3, 38, 54, 8, -28, -28, -15, -29, 14, 27, -43, 38, 3, -79, 89, 97, -100, -71, -1, 90, -5, -69, 78, 32, -18, 0, -8, -89, 54, 61, -80, 56, 9, -115, 64, 72, -53, 29, 43, -17, -58, 21, 18, -54, -32, -4, 42, -45, 17, 22, 46, 8, -25, 30, -48, -21, 8, 31, 1, -46, -19, 55, -10, -26, 49, 48, -44, -93, 99, -4, -110, 44, -3, 0, 81, -58, 20, 9, -82, 35, 31, -37, 46, 7, -5, -3, -13, 3, 29, -12, -43, 13, 17, 55, -14, -17, -5, 48, -1, -14, -68, 21, 5, -68, 23, 60, 8, -89, 73, 35, -54, -4, 22, -10, 0, 15, -11, -13, 20, 17, -27, -23, 27, 11, -79, 12, 81, 27, -47, -7, 8, -4, -5, -4, 38, 12, -30, -65, 59, 17, -26, 4, 11, -2, -7, 12, 12, -19, -1, 34, -2, -29, 9, 23, -19, -45, -73, 63, 68, -9, -55, -9, -13, 26, 74, 25, -47, -49, -17, -11, 60, 44, -6, -15, -51, 6, -3, -60, 102, -26, -23, 99, -59, 7, 12, -78, 49, 29, -14, 28, -70, -47, -2, 3, 90, -38, -56, 40, 0, 14, 29, -26, -28, 23, 41, 30, -78, -74, 107, -3, -98, 86, 70, -23, -20, -27, 30, 29, -111, 40, 38, -90, 82, 12, -59, 60, -29, 17, -32, -3, 30, -3, -30, 0, 19, 10, 34, -85, 74, 4, -65, -4, -22, 6, 61, 48, -22, 5, -34, 0, 21, -18, 44, -9, -94, 4, 27, -8, 0, -2, -12, 28, -6, -43, 29, 12, -30, 39, 60, -69, -41, -6, 17, 25, -1, -10, -12, -22, 82, 41, -24, 15, -68, 40, -17, -49, 25, -8, 55, 4, -12, 64, -80, 0, 21, -49, 13, -10, -9, 52, 35, -72, 47, 48, -25, -41, -74, 68, 43, -103, 22, 18, 0, 70, -74, 6, 17, -47, 0, 49, 66, -13, 26, -106, 9, 21, -43, 4, -9, 82, -59, -62, 10, 78, 76, -15, -53, -89, 53, 77, -77, -54, 95, 55, -99, -68, 62, 7, -26, 64, -30, -51, 72, -29, -43, 63, -26, 25, 41, -10, -2, -15, 35, 3, -27, 21, -9, 4, 45, -68, -4, -34, -11, 70, 1, 0, 2, -45, 26, -3, -93, -1, 32, 72, -53, 11, 20, -57, 36, 61, -47, -79, 48, 75, 36, -93, 8, 45, -88, 34, 69, -3, 1, -31, -26, 24, -31, -47, 93, -23, -73, 115, -49, -13, 72, -82, 0, 69, -6, -77, 21, 55, -46, -41, 42, -12, -22, 32, 11, 23, -47, -9, 43, -68, 48, 105, -43, -72, -30, 49, -9, 9, 30, -37, 17, -30, 12, 12, -71, 7, 25, 43, 44, -20, 22, -26, -9, -2, 1, 21, -89, -41, 102, 41, -111, 64, 30, -19, -30, 1, 30, -40, 13, 37, 55, -83, -80, 69, 18, -60, 55, 65, -108, 7, 63, -86, -17, 28, 27, -34, 30, 48, -77, 23, 89, -56, -25, 31, -77, 56, 10, -44, 15, 21, 17, -63, 52, 24, 8, -40, -12, 62, 0, 13, -40, -45, 39, 28, -12, -45, 15, 18, -21, 73, -72, -19, 12, 13, -10, -60, 72, -23, 9, 62, 21, -64, -90, 72, 70, -104, 34, 56, -40, 56, -44, -60, 9, -4, -29, -24, 41, 75, -6, -64, 37, 28, 23, -58, -43, 9, -7, 4, -8, 2, 68, 11, -64, 1, -28, 4, 9, -15, 62, -9, -72, 20, 17, 29, -2, -8, 1, 60, -45, 17, -8, -10, 73, -119, 43, 115, -107, -74, 122, -6, -72, 79, 2, -2, -54, -22, 114, -68, -13, 64, -78, 26, 61, -39, -34, -53, 63, 76, -105, -71, 91, -1, -80, 29, -7, 75, 11, -91, 23, -1, 13, 60, -32, -70, 57, 0, 22, 37, -45, 28, -32, 9, 53, -81, -3, -6, -22, 38, 51, -12, -31, 30, -14, 0, 37, -1, -14, -62, 17, 96, -64, -56, 46, 12, -14, -30, 37, 4, 5, 13, -80, 0, 1, 63, 7, -21, 56, 6, -75, 17, -8, 4, 26, -26, 26, -49, -4, -12, 0, 15, -49, 51, 47, -3, -24, -81, 102, -12, -75, 109, -23, -17, -26, 1, 41, -21, 3, -12, -13, 41, -18, -22, 44, 5, -23, -60, 69, 60, -70, -42, 73, 13, -105, 34, 8, -43, 66, -21, -32, 13, -47, 57, 85, -74, -28, 13, 14, 61, 2, -85, -8, 91, 1, -72, -11, 89, -22, -53, 39, 13, 14, 4, -85, 42, 13, -71, 2, 58, 17, -31, -37, -6, 23, 24, 30, -7, -52, -40, 54, 37, -13, -65, 19, 97, -27, -102, 76, 57, -44, 4, -18, -7, -14, 11, 14, -21, 55, 12, -54, -15, -17, -1, 64, 6, -66, 8, -2, -28, 57, 51, -77, -70, 94, 52, -81, -45, 85, -29, 13, 40, -28, 19, -81, -19, 8, 21, 72, -48, -49, 17, 23, 22, 15, 2, -83, 61, 95, -86, -54, 63, -36, -43, 82, 62, -103, 22, 12, -20, 15, -86, 22, 78, 22, -57, -52, 31, 77, -5, 6, -85, 34, 26, -62, 52, 3, -10, 1, -7, 12, 57, -78, 2, 10, 3, 64, -93, 26, 77, -89, -92, 108, 19, -11, 20, -38, 68, -63, -46, 61, 30, -19, -17, -30, -58, 12, 64, 20, 13, -34, -56, 70, 0, -76, 81, 5, -13, 9, -78, 64, 8, -55, 35, 51, -46, -57, 37, -3, -28, 80, 57, -88, -28, 42, -29, 2, 54, -55, -68, 69, 0, -9, 4, 1, 48, -49, 30, 30, -41, -22, -37, 80, 7, 2, 20, -19, -32, -78, 91, 48, -108, 40, 69, -28, -28, -48, -3, 2, -12, 19, 51, -8, 10, 54, 10, -32, -87, 64, -26, -15, 19, -60, 64, 23, -36, -26, 6, 17, 7, -10, -46, 32, 4, 26, 7, -46, 90, -21, -20, -35, 22, 28, -47, 54, -31, -11, -4, -4, 31, -27, -19, 28, 22, 46, -59, 7, 18, -53, 28, 3, 47, -19, -53, -37, 8, 42, 24, -11, -65, 3, 42, 45, 30, -93, 10, 0, -14, 94, -5, -73, -24, -22, 41, 109, -87, -106, 117, 19, -45, 34, -65, 23, -7, -27, 76, 1, -73, -8, 102, -52, -5, 54, -94, 25, 47, 4, 25, -56, 8, 19, -18, -37, -2, 48, -62, 22, 55, -80, 66, 6, -45, 0, 10, 58, -29, 0, -51, 7, 100, -86, -20, 95, -55, 18, 4, -95, 45, 6, -37, 35, 6, 56, -4, -82, -7, 42, 28, 23, -12, 4, -58, -58, 94, 40, 0, -24, -52, -29, -18, 28, -24, 76, -11, -56, 95, -29, -13, 6, -20, 56, 39, -103, 22, 31, -74, -4, 54, 89, -94, -45, 93, -68, 7, 53, -4, 29, -82, -55, 90, -9, -48, 90, -46, -38, 31, 24, 65, -97, -55, 43, 72, -39, -57, 98, -32, 1, -19, -64, 91, -29, 1, 49, -73, 30, -12, -53, 39, -6, 6, -1, -14, 90, -49, -36, 47, -18, 13, -20, 0, 44, 25, -40, 23, -10, -56, 14, -31, 15, 41, 36, 9, -48, -6, -40, -40, 74, 0, -21, 70, 3, -5, -32, -19, 76, -72, -81, 60, 27, 11, -52, -15, 35, 20, -12, 23, -32, -18, 105, -21, -65, 52, -13, -1, 21, -53, -18, -39, 58, 70, -79, -26, 63, -4, -43, 8, 32, -13, -39, -47, 108, -6, -59, 35, 8, 60, -75, -1, 61, -83, -20, 85, 57, -34, -6, -9, -88, 65, 41, -27, 24, -19, -34, -24, -22, 10, 77, -6, -1, 32, -31, -3, 24, 38, -85, -52, 98, -51, -52, 26, -21, 35, 0, -49, 0, 82, 26, -82, 37, 89, -90, -51, 70, -35, 17, 26, -2, 1, -71, 19, 9, 6, 13, -74, 49, 17, -13, 14, -28, 44, 17, -24, -31, 18, 31, -29, -6, 57, 18, -82, 35, 38, -20, -27, 26, -6, 0, 24, -5, -48, -69, 5, 48, 36, -69, -10, 56, 29, -20, 48, -19, -90, 22, 38, 20, 31, 31, -78, -1, 46, -51, 35, -26, -49, 7, -23, 58, -13, 4, 52, -87, 52, 34, -13, -26, -10, -26, 29, 17, -46, 80, -26, -2, -11, -76, 40, -3, 43, 74, -114, 2, 21, 9, 65, -27, -72, -47, 31, 2, 47, 64, -62, 6, 9, -75, 69, 88, -104, 9, -8, -17, 65, -30, -15, 30, 6, -1, 48, -42, -18, -42, -62, 94, 77, -108, -40, 119, -70, -5, 8, 0, 55, -52, 8, 39, 4, -34, 14, 36, -46, 6, 40, -96, 0, -1, 45, 6, -111, 97, 53, -36, 31, 12, -31, -5, 36, -71, -18, 79, 9, -9, -7, -27, -42, 2, -10, 73, -30, -104, 108, 28, -93, 18, 47, -6, 19, -14, -2, 39, -31, -39, 22, -2, -25, -8, -4, -8, 7, 88, -40, -72, 78, 39, 11, -77, -45, 24, -26, 13, 10, 61, 45, -61, -11, 1, -45, -15, 75, 62, -89, -42, 24, 22, 46, -20, 14, 37, -8, -66, 12, 60, -26, -19, 11, -19, 14, -51, -12, 98, -40, -90, 72, 1, -40, 41, -18, 23, 22, -29, -23, 44, 13, 2, -21, -32, 0, -7, 7, -30, 36, 22, -81, 9, 92, 21, -5, -4, -11, 0, -15, -52, 20, 32, -47, -18, 51, 47, 4, -18, -73, 4, 2, 52, -15, -15, 19, -13, -22, 5, 64, 14, -85, 4, 23, 3, 49, -95, 23, 12, 17, -15, -36, 42, -4, 26, 23, -43, -14, 28, 23, 22, -78, -58, 72, 14, -72, -39, 115, -7, -34, 93, -108, 14, 73, -85, 44, -11, -43, 43, 2, -26, 27, -31, 17, 21, -5, 41, -24, 1, -44, 24, 0, -34, 79, -57, -15, 116, -100, 10, -5, 0, 80, -114, 39, 19, -63, 61, -15, 27, -29, 9, 0, -4, 0, -94, 19, 83, 36, -3, -5, -99, 20, 82, -19, -35, 46, -12, -56, 82, -24, -60, 83, 29, -40, 9, -41, -79, 48, 31, 37, 20, -45, -51, 12, 43, -55, 35, 14, 1, 29, -13, 36, -64, -15, 13, 11, 6, 0, -19, -21, -25, 29, 40, 4, 12, -60, -35, 21, 78, -1, -28, 6, -52, 31, -1, -6, 0, -78, 9, 89, 63, -116, 38, -2, -21, 29, 7, 7, -80, -10, 75, -15, 20, 26, -102, 34, 51, -25, -53, 19, 80, 28, -85, -58, 61, 3, 27, 37, -52, -54, 36, 9, -58, 52, 6, -80, 82, 15, -71, 1, 6, 2, -15, 30, 7, -5, 63, -53, -8, 9, -32, 74, 14, -5, 14, -12, -94, 65, 0, -32, -8, 17, 87, -70, -15, -18, -15, 41, -20, 25, 20, -11, 25, 24, -73, -56, 17, 82, -18, 8, -20, -26, 81, -7, -10, -13, -20, 5, 27, -18, -26, 13, 22, -52, -31, -17, 21, 43, 3, 20, -23, -64, 9, 92, 47, -62, -52, -23, 15, 41, -37, 0, 12, 44, -7, 1, 29, -31, 29, -57, -24, -17, 49, 89, -91, 20, 70, -51, -27, -15, -28, 38, 5, -17, 44, -58, 32, 77, -83, -37, 6, -6, 48, 22, -75, 62, 21, -47, 56, -81, 9, 119, -99, -27, 93, -59, -6, 28, 25, -59, 13, -1, -20, 19, -20, 24, -40, 36, -31, -9, 89, -44, 5, 25, -24, 61, -25, -91, 37, 4, -61, 48, -9, -23, -1, 63, 27, -9, 5, -60, 64, -5, -60, 43, 13, -77, 46, 83, -41, -76, -17, 45, -9, -34, 72, -11, -82, 47, -13, 44, 28, -49, -17, 20, 36, -20, -6, -26, -30, 87, 26, -76, -29, 77, 55, -13, -88, 12, 66, -42, 48, -61, -85, 39, -5, 79, 7, -63, 10, 14, -18, 19, 77, -38, -49, 22, -58, 32, 86, -90, 31, -2, -34, 0, -34, 25, 73, -11, -74, 51, -31, -46, 81, -25, -27, 99, -61, 3, 34, -53, 15, 13, -8, -17, -22, 28, 95, -80, -24, 65, -35, -17, 65, -68, -15, 29, -42, 59, -7, 21, -25, -17, -23, 32, 68, -51, 22, 23, -28, -57, -3, -32, 47, 75, -51, -63, 15, 41, -36, -6, -22, 41, 88, -93, -1, 70, -66, -18, -5, 60, -22, -28, 43, -47, 28, -25, 37, 26, 0, 6, -29, -1, -28, 40, -58, 35, 61, -40, -31, 27, 63, -59, -18, 37, -22, -18, -22, 24, 48, -25, -25, 48, -57, 14, 1, -48, 103, 36, -112, 13, 40, -30, -7, 13, 9, -65, 49, 47, 27, -98, -9, 88, -46, -23, -6, 43, 42, -28, -20, 0, -36, -46, 30, -1, 61, 9, -29, 76, -69, -6, 66, -29, -14, -52, -12, 80, -5, -73, 41, 18, -62, 34, -23, 3, 95, -29, -41, 47, -40, -62, 28, 15, -18, 35, 37, -47, -48, 31, 2, -6, 24, -38, -32, 97, -1, -44, 70, -11, 11, -1, -81, -28, 9, -14, 66, 83, -22, -63, 19, 47, -17, -61, -46, 75, 62, -5, -87, 35, 24, -82, 29, 26, -10, -3, 12, 5, -27, -29, 18, -38, 60, 26, -86, 72, 9, 2, 63, -105, -39, 62, 32, 29, 1, -102, 17, 62, -20, 42, -13, -86, -18, -4, 31, 58, -8, -39, -47, 75, 19, -53, 62, -35, -5, -3, -74, 6, 86, 80, -96, -45, 49, -43, -13, 29, -30, -17, 70, 81, -86, -53, 107, -18, -55, 27, 61, -65, -9, 11, 8, 8, -39, 70, -27, -42, 43, 9, -36, 42, -24, 0, -23, 5, 66, -35, -74, 34, 56, -4, 6, -9, -38, 0, -28, 17, 31, -98, 65, 108, -86, -11, 1, 7, 34, -25, -11, -32, -15, 63, -13, -40, 65, -38, -12, -2, 38, 22, -78, 6, 14, 38, -23, -19, 38, -52, -1, 46, -14, -48, 44, 9, 25, 45, -70, -29, 20, 8, 23, 3, -37, 31, -36, 5, 108, -51, -85, 34, 80, -55, -68, 8, -15, -3, 80, 0, -30, -32, 47, 61, -82, -18, 93, -39, -83, 26, 20, 24, 34, -44, -60, -2, 78, -7, 4, 72, -38, -59, -5, 45, -24, 15, 34, -40, 36, 0, -19, 3, -34, 51, -70, 18, 34, -110, 93, 36, -81, 2, 81, -46, -42, 21, -49, 34, 12, -20, -27, 88, 5, -29, 23, 1, 5, -55, -15, 17, 59, -56, 23, 26, -27, 89, -91, 4, 112, -111, -45, 27, 2, 18, -41, 73, 14, -65, -3, 26, 22, -31, 4, 47, -41, -83, 52, 52, -46, 17, 72, 8, -20, 4, -56, -25, 69, -37, -17, 46, -11, -86, 54, 104, -71, -74, 64, 55, -29, -53, -5, -9, 24, 1, -94, 97, 5, -40, 38, -21, -3, -2, 10, -23, -20, 43, 62, -63, -78, 44, 73, 0, -41, 39, -10, 19, -36, -56, 74, 20, 6, -65, 32, 31, -87, 77, -8, -56, 37, 4, 36, 32, -89, -44, 10, -18, 91, 51, -58, -81, 6, 13, 7, 56, 52, -92, -12, 12, -36, 40, 35, -30, -24, 73, -23, 23, 11, -10, -10, -63, 15, 22, -51, 21, 69, -62, 25, 69, -100, -34, 78, -3, -21, 0, -36, 29, -2, 40, 20, -17, -12, -35, -26, -37, 13, 64, -36, 27, 52, -47, -9, -65, 89, 24, -41, 47, -18, 3, -19, 17, -31, -52, 15, 37, 36, -19, -43, 55, 19, -23, 37, 6, -56, -10, 80, -41, -60, 68, -15, -7, 22, -52, 62, -25, -3, 39, -93, 4, 20, 0, 1, -30, 59, 14, -80, -15, 105, -13, -74, 34, -15, -36, 20, 19, 65, -31, 0, 23, -77, 8, -5, 31, 68, -55, -79, 65, 70, -61, -40, -18, 48, 48, -47, 21, -47, -14, 93, 34, -6, -69, -43, 89, -19, -22, 19, -46, -32, -2, 71, -19, -13, 62, 32, -36, -85, -25, 7, 79, 5, -55, 85, -39, -96, 38, 71, -56, 21, 77, -111, 14, 92, -42, -4, -15, -44, -8, 28, 11, -9, -11, 12, -3, -60, 48, 48, -53, 5, 57, 23, 30, -89, -2, 104, -77, -74, 62, -1, -51, 7, 0, 75, -34, -18, 71, -72, 48, 37, -20, -28, -81, 77, 73, -107, 42, 7, -37, -11, 13, 19, 10, 44, -70, 31, 9, -12, -42, -58, 102, -5, -52, 12, -42, 25, 82, 5, -22, 39, -46, -20, -14, -15, 38, 37, 8, -35, -40, -27, 41, 61, -8, -32, -7, 51, -3, -108, 39, 42, -51, 7, 38, 7, -3, 19, -57, -11, 22, 31, 5, -22, 8, -6, -37, 44, 27, -26, 9, -14, -32, -61, 47, 48, -4, 41, -11, 11, -45, -82, 56, -8, 17, 73, 22, -75, -21, 75, 23, -110, 19, 25, -20, 9, -5, 75, -58, -62, 46, 40, 13, -8, 2, -28, -52, 20, -10, 48, 8, -53, -30, 42, 49, -14, 25, -20, -71, 3, 36, 42, 5, -57, -19, -18, 62, -22, -54, 4, 4, 82, 45, -70, -14, 45, 9, -69, -43, 2, 69, 54, -51, -52, 7, -3, 44, 11, -22, -27, 17, 12, 12, 23, -43, -3, 3, 18, -47, 65, 0, -21, 56, -45, -72, 38, -21, 32, 59, -65, -52, 15, 102, -17, -32, -2, 0, 9, 9, -21, -15, 25, -8, 0, 48, -55, -3, 54, -39, -26, -17, 93, -49, -71, 49, -30, 57, 28, -87, 5, 72, -30, -86, 65, 61, -10, -49, -24, 0, 48, 41, -14, -11, -60, 5, 12, -1, -18, 46, 72, -48, -57, 55, 9, -15, -29, 2, 40, -25, 51, -69, -39, 18, -43, 3, 58, 60, -43, -79, 81, 3, -36, 66, -32, 38, -64, 5, 34, -86, 77, -29, 3, -5, 25, 14, -23, -3, 17, 17, -28, 68, -49, -66, 64, 18, -65, 37, -35, 0, 46, 24, 27, -81, 0, 15, -69, 51, 3, -54, 80, 54, -59, -29, 70, -35, -14, 48, -42, 23, -47, -46, 71, -7, 0, 2, 10, 44, 14, 0, -44, -29, 47, -41, 1, 26, -47, 70, -56, -19, 12, 22, 34, -48, 17, -31, 48, 0, -95, 30, 0, -51, 77, 47, -37, -14, -41, -4, 27, -22, -26, 75, 36, 19, -54, -52, 45, 10, -4, -8, -9, 8, 13, 24, -40, 28, 14, -102, 28, 9, 20, 7, -14, -13, 56, 55, -30, -73, -61, 110, -9, -88, 75, 49, -70, 19, -1, -24, 29, -5, -31, 19, 2, -18, 43, -37, 10, 37, -25, 17, 72, -96, -65, 53, -1, -7, 0, -30, 8, 28, 58, 1, -37, 43, -64, 27, 38, -64, 5, 45, 42, -29, -23, -46, -24, 0, 5, 79, 14, 3, 5, -28, 38, -62, -82, 38, 17, 8, -11, 27, 57, -46, -63, 43, -27, -15, 52, -8, 29, 56, -51, -19, 49, -98, 23, 113, -98, -55, 76, 49, -55, -30, 46, -40, -1, 54, -1, -70, -48, 95, 66, -104, -36, 1, 26, 25, -9, -31, 35, 39, -91, 7, -1, 46, 21, -88, 49, 34, -34, 17, -25, 22, 73, 20, -107, -15, 75, -19, 4, 23, -10, -40, 31, 38, -38, -25, -49, 62, 27, -9, -8, -40, -4, -9, 8, -5, 15, 36, 29, 2, -37, -89, 45, 13, 24, 28, -2, 10, -81, 22, 8, 19, -15, -66, 60, 32, -4, 11, 7, -66, 0, 87, -17, -1, -34, 12, -9, -22, 73, -93, 4, 9, -69, 31, 4, 66, 59, -88, -12, -21, 24, 90, -24, 28, -69, -52, 60, 35, -41, -42, -29, 71, 21, -45, 69, -14, -9, -55, -11, 38, -35, -25, 28, 9, -19, 55, -11, -71, 79, 62, -93, 14, 59, -96, 22, 79, -37, -25, 6, 30, 17, -23, 11, -52, -45, 59, 24, 34, 4, -75, -39, 80, -14, -7, -20, -11, 47, -59, 53, -4, 2, 91, -105, -23, -8, 28, 32, -43, 2, 38, 8, -94, 39, 0, -52, 82, 37, -5, 24, -49, -61, -13, 9, 15, 66, -11, -81, 3, 40, 56, -2, -43, 32, 26, -92, 27, 57, -59, -17, 59, -15, -28, 78, -3, -6, -64, -11, 49, -71, -6, 91, -42, -19, -9, -4, 46, -42, 27, 24, 20, -8, -69, 1, 2, 47, 20, -78, -3, 70, 11, -55, -37, 6, 0, 72, -20, -63, 61, 6, -22, 55, -11, -43, 32, -21, -45, 57, 47, -21, -5, -23, -28, 15, 66, -27, -23, -24, 2, 82, -66, -70, 26, -14, 29, 5, 60, 5, -36, 9, 31, -40, -47, 24, 4, 76, -19, -18, 42, -65, -18, 14, 1, 63, -81, -18, 37, -13, 44, 41, -41, 0, -28, -37, 98, -25, -10, 69, -110, -23, 55, 13, 25, 6, -51, -58, 81, 37, -77, 14, -26, 15, 7, -22, 80, -76, -14, -20, 43, 27, -91, 25, 5, -29, 100, -26, -31, 112, -96, -4, 62, -41, 31, -27, -8, -43, 27, 49, -5, -24, -71, 106, -34, -60, 83, 19, 1, -68, 23, 44, -63, 47, 44, -34, -71, 30, 70, -105, 10, 86, 0, -37, -43, 28, 47, -73, -13, 74, -21, -17, 24, 40, -26, -98, 2, 31, 36, -17, -34, 60, 23, -75, -2, 68, 0, -75, -9, 68, -69, 1, 43, -65, 54, 91, -38, 10, -74, -27, 60, 13, -43, -23, 57, 14, -9, -49, -40, 24, 19, 37, -24, -66, 75, 59, 2, -37, 4, 17, -103, 47, 105, -56, -109, 68, 32, -35, 56, -39, -41, 3, -22, 3, 71, 36, -69, -52, 98, -21, -27, 29, -94, 61, 48, -21, 31, -37, -37, 11, 68, -27, -47, 63, 26, -46, 18, -29, -58, 53, 18, 15, -76, 20, 17, -6, 57, -52, -35, 18, 60, -61, -82, 78, 87, -34, -30, 28, -74, 43, 17, -3, 17, -32, 81, -70, -54, 77, -10, -1, 17, -78, 14, 29, 31, 32, -66, 0, -22, 9, 0, 19, 60, -88, 10, 31, 10, -20, -74, 73, -1, -52, 69, 12, -60, 15, 55, -4, -18, -44, 17, -26, -9, 9, 6, 22, 39, -37, -89, 19, 60, 21, -71, 11, 43, 47, -66, -31, 24, -27, 22, 0, 52, -23, -72, -6, 81, 72, -12, -24, -61, 2, 39, 19, 10, -44, -46, 52, 7, -45, 74, -43, -3, 0, -31, 41, 24, 13, 10, -61, 6, 28, -60, 62, -14, -22, 52, -21, -42, 61, -72, 8, 42, -30, 49, -61, -49, -19, 82, 45, -64, 45, 25, -70, 45, -6, -27, 72, 4, 5, -105, 35, 10, -51, 76, -3, -51, 14, -25, 17, 55, -93, 27, 72, 8, -31, -96, 69, 34, -10, 4, -10, 54, -85, -56, 75, 20, -82, 37, 26, 8, 44, -49, -68, 15, 2, 20, 56, -3, 17, -18, -40, -55, 10, 10, 43, 66, -86, 25, 8, -78, 26, 2, -43, 34, 37, 10, 54, -25, -42, -11, 6, -19, 27, 30, -25, 53, -40, -61, 71, -46, 34, 6, -99, 45, 15, -29, -22, 43, 86, -35, -10, 0, -31, 55, 31, -85, -24, 83, 0, -66, -36, 7, 1, 80, 40, -110, 21, 108, -63, -19, -24, -28, 76, -34, 18, -17, -63, 106, 21, -69, -17, 11, 19, 60, -45, -35, -26, 42, 25, -25, -21, -31, 95, -21, -38, 19, 0, -17, -3, 51, 48, -27, -62, 11, 71, -70, -4, 28, -76, 19, 48, -3, 32, -21, -34, -10, 29, 49, -80, -30, 23, -12, 51, -14, -10, 8, 3, -9, -10, 22, -71, 39, 82, -21, -58, 40, 40, -63, -62, 77, 43, -12, -15, -12, -36, 36, 88, -115, -21, 119, -59, 2, 15, -97, -13, 95, 1, -7, -24, -9, 124, -98, -55, 95, -10, -6, 24, -80, 40, 72, -114, -2, 56, -19, -36, 22, 19, 25, 40, -115, 36, 92, -1, -83, 19, 5, -103, 22, 83, -13, -96, 97, -1, -40, 57, 7, -24, -53, 63, -6, 0, 60, -10, -34, -51, -24, -35, 59, 92, -15, -31, 37, -14, -13, -45, -15, 82, -58, 6, 56, -74, 44, 17, -55, 22, -35, -43, 86, 22, -92, -5, 18, 78, -38, -13, 30, -85, 60, 88, -81, -44, 75, -46, -58, 40, -3, 39, -10, -37, 46, 20, 24, -22, -48, -30, 88, 4, -71, 64, 23, -31, -55, -44, 46, -4, 31, 56, -66, 4, 29, -18, -41, -25, 48, -7, -5, 46, 28, 3, -80, -14, 22, 32, 51, -25, -83, 28, 88, -45, -15, 2, 31, 14, -40, -29, 30, -8, 5, 74, -5, -51, -56, 66, 6, -7, -30, -88, 41, 87, 3, -37, -39, 47, 15, -100, 22, 18, 42, -21, -3, 23, -19, 29, 39, -59, 0, 70, -72, 26, 31, -56, -28, -20, -9, 71, 63, -63, 6, 12, -68, 8, 62, 3, -53, -29, 15, 58, -8, -53, 58, -14, -28, 37, 15, 10, -27, 38, -31, -76, 66, -23, -19, 17, -65, 107, -25, -90, 43, 70, 10, -23, -9, -13, -19, 26, 44, -5, -4, -56, -37, 30, 19, 46, -44, -53, 54, 41, -37, 21, -12, -81, 0, 57, 24, -62, 57, -3, -22, -14, -19, -10, 48, 60, -45, 51, -6, -89, 46, 77, -56, 11, -2, -13, 54, -47, -44, -1, -5, 29, 0, -40, 59, -1, -69, -26, 47, 73, -26, -83, 56, 62, -95, 19, 6, -7, 49, -20, 36, -19, -30, 2, -31, 78, -12, -86, 34, 30, 0, 28, -49, 22, -12, 10, 23, -105, 99, 44, -6, -41, -17, 51, -5, 21, -44, -85, 12, 90, 6, -59, -17, -23, 29, 63, -76, 18, 88, -43, -41, -1, -15, 21, 0, -27, 34, -2, 1, 19, -44, -4, 65, 48, -68, -26, 72, -23, -1, -26, -20, 4, 2, 54, -20, -56, 5, 36, -41, -15, -4, 7, 71, -20, -78, 69, 61, -43, -23, -27, -23, 20, 54, 44, -40, 7, 36, -83, 8, 10, 4, -32, 17, 6, 20, -1, -49, 27, 12, 22, -13, 30, -59, -34, 6, -25, 15, 48, 43, -30, 22, 15, 11, -13, -30, -6, -7, -17, 22, -20, -3, 25, -54, 13, 34, -31, -8, 96, -8, -83, 30, -23, 34, 63, -75, 43, 34, -40, 0, -13, -48, 18, 3, -34, -14, 63, 45, -22, -41, -44, 70, 44, -38, 35, -31, -94, 0, 70, -18, -25, 100, -11, -27, 42, -41, -85, 86, -28, -9, 64, -41, -35, -49, 74, 15, -61, 29, 60, 25, -12, -73, 4, 30, 0, 21, -21, 15, 23, -62, 17, 15, -75, 7, 79, 57, -31, -92, 30, 49, 5, -12, -102, 81, 24, -24, -13, -17, 24, -64, 10, 98, -25, -92, 18, 83, 17, -3, 9, -48, -43, 4, 58, -28, 13, 47, -62, -21, 66, -30, -81, 75, 42, -74, 46, -21, -77, 9, 53, 37, -55, -22, 24, 29, -27, 42, 24, -102, 60, 10, -35, -6, 15, 24, -37, 55, -64, 34, 8, 5, 2, -74, 86, 21, -10, -3, 0, 21, 4, -36, -29, -51, 30, 82, -21, -85, 36, 1, -74, 77, -8, 2, 47, 31, -66, -80, 85, -18, -70, 95, -10, -66, 21, 71, -22, -100, 69, 64, 31, -37, -57, 0, 20, -26, -26, 3, -22, 102, -18, -73, 64, -5, -49, -1, 25, -24, 9, 90, -43, -37, 76, -55, 5, 98, -94, -15, 106, -26, -41, 48, -68, 13, 24, -46, -8, -22, 68, -32, -30, 48, 6, 10, 43, -21, -81, -42, 64, 18, 26, 42, -108, -8, 96, 9, -45, 24, 13, -54, 18, -25, -27, 64, -34, 0, 18, -43, -20, 64, 35, -54, 24, -47, -22, 44, 22, -13, 6, -25, 24, 55, -120, 53, 21, -19, 62, -24, 28, -37, -55, 24, 25, 26, -21, -95, 26, 88, -49, 7, 39, 5, -26, -46, -38, 40, 87, -17, -61, -20, 89, -36, -98, 106, -6, -75, 86, 54, -80, 4, 18, -26, 27, -65, 2, 94, -47, -80, 69, 32, -74, -1, 41, -10, 40, 2, -60, 38, -15, -10, 20, -60, 64, 30, -63, -53, 87, 21, -111, 30, 0, 20, -14, 8, 66, -12, -6, 15, 38, -52, -37, -35, 35, 95, -45, -9, -14, 26, 3, -28, 18, 0, 44, -29, -56, -21, 26, 10, -19, 29, 15, 3, -62, 22, 10, 4, 7, 1, 44, -66, -26, -15, 8, 10, -51, 75, 88, -64, 12, -1, -74, 28, -1, -26, -22, 32, 43, -17, 44, 46, -78, -30, 47, -28, -29, 60, -23, -19, 60, 17, -62, -78, 2, 37, 22, -49, 27, -4, 17, 18, -24, 57, 20, 0, -82, 19, 31, -41, 26, -36, 6, 36, 45, -58, -80, 15, 91, -14, -1, 62, -89, -63, 76, 5, -47, 99, -45, 1, -18, -5, 17, -41, 51, 36, -41, -31, 57, -11, -47, -48, 64, 43, -10, 2, -14, 17, 20, -35, 23, 39, -87, -62, 64, 77, -55, -71, 63, 34, -95, 48, 28, -79, 9, 56, 68, -32, -61, 14, 65, -24, -34, 41, -73, -21, 19, 24, -27, 41, 10, -116, 83, 10, -62, 14, 92, -7, -57, 46, 23, -18, -37, 54, 10, -29, 22, -11, -45, -41, 7, 0, 24, 65, 19, -26, -47, -48, 0, 12, 83, -11, -77, 53, 1, -30, 69, -17, -20, 32, -83, 26, -8, -8, 57, 3, -15, -31, -5, 26, 18, -19, 49, -49, -44, 71, 13, -2, 0, 35, -80, -5, 22, -46, 26, 0, 59, -40, 6, 37, -30, 58, -71, -14, 47, -13, -13, 30, -45, -18, 57, -30, -13, -25, 34, 28, 42, -42, -62, 63, -31, -27, 36, -29, 38, 39, -4, -17, 19, 21, -93, 12, 55, -52, 0, -29, 48, 71, 0, -85, -36, 57, -25, 39, 30, -82, -19, 73, -38, 31, 3, -43, 2, 14, 59, -72, -31, 51, 19, -8, -59, 63, -21, -2, 12, -45, 104, -53, -62, 100, -27, -96, 26, 56, 56, -76, -1, 35, -5, -18, -44, 0, 26, 47, 18, -25, -4, 6, -85, 18, 83, -29, -52, 88, -36, -42, 65, -69, 40, 0, -77, 12, -5, 39, 70, -60, -13, 65, -24, -17, 24, 42, -20, -37, 0, 17, -62, -24, 115, -56, -3, 88, -68, -34, 38, 30, -76, -26, 76, 53, -46, 22, -49, -29, 62, -4, 43, -65, -26, 15, 25, 0, -52, 7, 49, 61, -109, 11, 34, 4, -23, -80, 94, -2, -1, 22, -81, 32, 83, -5, -3, -54, 13, 55, -82, -34, 75, -64, 13, 27, -47, 41, 2, 35, -64, -35, 94, -64, -21, -2, 56, 42, -79, 37, 59, -60, -54, -1, -27, 10, 86, 58, -43, 10, 0, 5, -23, -56, 76, -35, -27, 29, 3, -2, -68, 55, 52, 1, 12, -59, -88, 68, 70, -56, -5, 20, -4, 27, -2, -9, -53, -5, 45, 11, 5, -63, 19, 70, -9, -14, -55, -13, -4, 39, 72, -74, 5, 32, -48, -4, 63, -25, -46, 21, 49, -53, -66, 44, 61, 43, -77, -79, 36, 60, 25, 17, 19, -43, -6, 28, -59, -59, -5, 25, 72, 45, -26, -13, -12, -56, -15, 30, 8, 25, 54, -52, -5, -14, -7, 57, 5, 28, -23, -48, -2, 21, -35, 15, -22, -38, 24, 7, -4, -3, 55, -23, -45, 29, 52, 28, -28, -54, -28, -21, 83, 3, -72, 76, -12, -57, 20, 13, -28, -22, 57, 59, 0, -66, -38, 88, -17, -9, -14, 0, -13, 18, 90, -63, -42, 48, -13, -70, -24, 48, 0, 37, 53, -48, 3, 37, 24, -88, -58, 107, 0, -114, 76, -3, -68, 18, 64, 26, 5, -39, -65, 11, -19, 2, 40, 29, 30, 28, -42, 26, -36, -19, 63, 14, -46, -46, 76, -45, -21, 20, -73, 91, -3, -14, 87, -53, -87, 59, -5, -102, 113, 17, -87, -18, 18, 62, 10, -40, 0, -7, -35, 53, 83, -82, -18, 34, -18, 36, -9, -37, 30, 53, -59, -62, 59, 4, -26, 88, -70, -9, 5, -69, 9, 6, 5, 8, 73, 12, -8, -37, 0, 89, -97, -2, 3, -4, 7, -11, 31, -4, -25, -47, 49, 0, 3, -25, 26, 0, -72, 72, 80, -87, 4, 89, -80, 29, 5, -97, 43, 82, -23, -62, 59, 12, -92, 63, 9, -82, 53, 19, 27, 0, -2, -37, 23, 0, -63, 53, -25, 0, 12, -59, 46, -4, 6, 99, -88, -73, 0, 68, -12, -21, 6, 23, 102, -86, 1, -2, -34, 29, 18, 13, -79, 14, 88, -78, 15, 26, -25, -8, 26, -12, -68, 73, -20, -37, 38, 7, -22, 38, -37, -13, 13, -30, 35, -19, 17, 11, -18, -17, 42, 0, -25, 74, 17, -47, 14, 32, -24, 11, -88, 2, 87, -41, -55, 70, 30, -21, -11, -80, 15, 39, -2, 12, 9, 29, 11, -64, -46, -6, 6, 86, -26, 4, 66, -103, -20, 59, 42, -43, -58, 66, 68, -85, -65, 34, -39, 79, -7, -73, 114, -12, -9, 19, -95, 21, 26, 8, 51, -42, 22, -34, -47, 17, -29, 0, 7, 37, 61, -60, 12, 20, -107, 83, 24, -57, -18, 10, 22, -51, 76, 0, -41, 64, -4, 0, -49, 46, 6, -2, 25, -79, -32, 68, 26, -85, 69, 34, -24, 15, -3, -11, 13, 22, -44, -47, -32, 25, 54, -30, 0, 13, -9, -20, -32, -11, 66, 28, -77, -13, 25, 37, -3, -3, -3, 20, 42, -48, -31, 14, 76, -37, -106, 93, 73, -36, -89, 66, -12, -37, 36, -11, -20, 3, 79, -78, 14, 36, -48, 49, -3, 1, -25, 13, -4, -31, 37, 14, 30, 2, -56, -4, 75, -53, -20, 41, 19, -2, -4, -82, -14, 9, -4, 53, 17, -35, -3, 29, -2, -30, -31, -3, 58, 52, -100, -32, 17, 44, -17, -59, 51, 13, 48, -7, -15, 49, -82, 25, 46, -108, 55, 8, -93, 53, 38, 34, 15, -53, -25, 11, 6, 29, 9, -20, -28, 18, 31, -6, -44, 13, 41, 3, -61, 0, 15, -78, 28, 26, 40, 53, -57, -15, 60, -19, -76, 12, 13, 28, 48, -10, -47, -37, 43, -60, 31, 104, -41, -24, 4, -65, -9, 24, 29, 22, 4, 45, -34, -58, -21, 26, -28, 32, 11, -77, 15, 23, 23, 31, -35, -17, 19, 3, 60, -70, -32, 90, 30, -53, -46, 39, -27, 31, 64, -88, -37, 90, -45, -71, 11, 23, 46, -12, -52, 56, 15, -35, -29, 64, -7, -66, 47, 10, -39, -26, 52, 37, -48, -3, -15, 17, 12, -42, 51, 54, 4, -99, 32, 71, -82, 48, -17, -12, 31, -68, 44, 24, 7, 15, -20, 19, -31, -86, 32, 20, -20, 63, 57, -46, -31, -49, -29, 72, -2, 22, 11, 21, -55, -64, 92, -24, -40, 77, -38, -9, 8, 4, 38, -98, 42, 15, -96, 104, 19, -62, 9, 21, 22, -45, -24, 80, -4, -53, 40, 12, -8, -57, 37, 20, -9, -5, 17, -26, -60, 92, 49, -52, 9, -24, -13, 29, -29, 23, -3, 13, -40, 7, 32, -18, -38, 8, 64, -45, -22, -6, -29, 56, 23, 5, -11, -74, 1, 94, -11, -59, 99, -54, -89, 88, 9, 8, -17, 3, 31, -22, 15, -8, 6, -61, -24, 58, 36, 38, -75, -74, 31, -17, 70, 56, -97, -52, 90, 12, -65, -34, 87, 7, -85, 0, 69, 59, -104, -35, 60, 36, -57, -30, 28, 40, -3, 2, 7, -54, 41, 20, -37, 51, 26, -57, -4, 40, -1, -22, -54, 40, 53, -77, -61, 81, 10, 9, 28, -74, -2, -44, 76, 26, -75, -2, 68, 29, 0, -35, -4, 40, -14, -20, -19, 11, 30, -23, -59, 32, 42, -1, -36, -13, 29, 11, -44, -45, 21, 73, -25, -4, 48, -40, -65, -26, 43, 92, 5, -44, -37, 22, -4, -51, -18, 69, 49, 12, -44, -96, 44, 86, -8, 8, -18, -68, 21, 26, -24, 43, -11, -27, 40, 15, 44, -48, 10, -3, -48, 40, -72, 27, 41, -98, 91, 20, -121, 51, 35, -76, 44, 58, 31, -57, -21, 12, -12, -22, 19, 97, -93, -78, 65, 57, -62, -1, 30, -49, -25, 72, 79, -96, 13, 5, -59, 80, 1, -42, -2, 38, 13, -74, 8, 44, -18, -35, 38, 80, -62, -28, 66, -43, 1, 22, -97, 49, 108, -65, -90, -5, 6, 78, -8, 0, 82, -48, -11, -4, -71, -14, 10, 32, 1, 21, -28, -15, 94, 5, -24, -57, 0, 14, 10, -17, 17, 48, -80, 14, 94, -82, 10, 11, -97, 20, 12, -35, 61, 94, -62, 14, -35, -27, 47, -32, -6, 13, -26, -23, 23, 38, 6, 24, -34, -72, 6, 73, 66, -73, 0, 48, -25, 11, -71, -7, 122, -81, -20, 92, -77, -60, 85, -23, 25, 0, -31, 17, -7, 54, -8, -74, 0, 20, -71, 58, 39, -65, 41, -8, -3, 19, 39, -6, -83, -8, -14, 18, 0, 78, -24, -54, 18, 37, 56, -70, -52, 22, 36, 52, -36, -59, -20, 53, 51, -89, 0, 87, -19, -92, 80, 85, -76, 34, -35, -26, 1, -71, 105, 2, -102, 82, 56, -87, 31, 1, -42, 68, 23, -94, 10, 98, -68, -5, 41, -19, 34, -73, -18, 12, -53, 41, 76, 5, -38, -46, -19, 51, -3, -46, 52, 27, -76, -1, 55, 41, 0, -77, 20, 20, -62, 35, -13, 5, 2, 29, -9, 13, 68, -28, -83, 38, 9, -6, 43, -28, -53, 22, 23, -76, 91, 49, -26, -77, -39, 29, 54, 47, -48, -10, -42, 0, 110, -57, -80, 0, 83, 19, -96, 40, 98, -69, -32, 17, -54, -10, 80, -13, -7, 104, -71, -8, 65, -98, 1, 114, -68, -30, 48, 15, -68, 6, 42, -92, 63, 48, -92, 36, 64, -55, -31, 49, 10, -86, 46, 70, -98, 15, 75, -86, 8, 1, 17, 54, -96, 42, 31, -30, 9, -28, -13, 52, -40, 5, 94, -92, -36, 24, -54, 9, 58, 24, -47, -41, 71, -24, 6, 86, -8, -8, -90, -2, 102, -71, -58, 7, 60, 61, -22, -17, -58, -15, 11, 11, -8, -25, 35, 44, -22, -14, 51, 56, -82, -88, 13, 76, 0, -92, 75, -8, -11, 76, -7, -19, 3, 42, -12, -23, 11, -14, -65, 47, 58, -53, -49, 49, 29, -12, -17, 25, -8, -76, 83, -4, -51, -11, -39, 60, -13, 15, 53, -6, 0, -46, -6, 1, -4, -19, -19, -11, 57, 3, 36, 4, -27, 6, -61, 27, -30, 35, 30, -39, -14, -19, 69, 21, -52, 55, -32, -44, 70, 17, -29, -41, -25, 53, 51, -49, 35, 30, -44, -1, -54, -6, 94, 5, 0, -54, -79, 82, 68, -45, -66, 52, 45, 0, -15, -96, 53, 39, -29, 10, -28, -60, 58, 32, -3, -1, 1, 49, -85, -19, 25, -26, -23, -10, 93, 63, -65, -74, 56, 1, -34, 99, -57, -73, 98, 11, -57, 40, -36, -65, 28, 22, -10, -43, 58, 93, -44, -26, 28, 0, -45, -75, 87, 18, -88, 94, -29, -43, 109, 3, -17, -12, -9, 55, -90, -19, 68, -37, 0, 11, 9, 29, -75, -1, 95, -17, 2, -41, -25, 30, -62, 19, 49, 5, 38, -15, -14, 27, -39, -19, 54, -61, -34, 46, -27, -10, 5, 21, 64, 3, -57, -15, 32, -21, -19, 15, -13, -39, 65, 51, -29, 26, -19, -72, 51, 15, -87, 36, 21, -12, 18, -56, 40, 68, -9, -76, -31, -5, 58, 8, 0, 1, -7, 31, -21, -24, 27, 76, -68, 3, 37, -76, 27, -4, -31, 59, -11, 13, -17, -77, -1, 88, -22, -70, 46, 79, -56, -7, 95, -92, -87, 95, 17, -93, -4, 109, -7, -86, 72, 56, -85, -3, 6, -78, 82, 62, -18, -19, -11, -35, -6, 80, 27, -6, -81, -13, 71, -28, -17, 34, -9, 6, -2, 9, 24, -8, 27, -75, -73, 77, 72, -45, -34, -34, 9, 23, 30, -6, 4, 17, -44, 20, -15, 7, -10, 12, -4, -49, -18, 88, -36, -24, 95, -43, 6, 7, -28, 11, 22, 9, -21, 4, -11, -80, 61, 88, -55, 3, -9, -31, 19, -54, -30, 94, 42, -40, 19, -76, 19, 115, -123, 7, 87, -28, -11, -22, 0, -41, -8, 20, -31, -27, 6, 44, 2, -40, 20, 80, -63, 13, 51, -44, -40, 20, 47, -2, 4, -68, 56, 24, -89, 69, 29, -115, 64, -6, -21, 41, -46, -27, 41, 36, -78, 48, 81, -78, 25, 13, -111, 96, 3, -57, 51, -39, -34, 76, 70, -31, -79, 38, -9, -56, 86, -2, -35, 13, 15, -56, 32, 82, -88, -13, 3, -31, 10, 64, 19, -51);
                                                      
    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project
 
    constant SCENARIO_ADDRESS : integer := 0;    -- This value may arbitrarily change
 
    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
 
                o_done : out std_logic;
 
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;
 
begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
 
                o_done => tb_done,
 
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );
 
    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;
 
    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data;
                    tb_i_mem_data <= tb_o_mem_data after 2 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 2 ns;
                end if;
            end if;
        end if;
    end process;
 
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
 
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;
 
        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
 
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;
 
        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';
 
        -- Wait some time for the component to reset...
        wait for 50 ns;
 
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
 
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock
 
 
        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        wait until falling_edge(tb_clk);
 
        memory_control <= '1';  -- Memory controlled by the component
 
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
 
        tb_start <= '1';
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        wait for 5 ns;
 
        tb_start <= '0';
 
        wait;
 
    end process;
 
    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin
 
        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';
 
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
 
        wait until rising_edge(tb_start);
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);
 
        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE 1)" severity failure;
    end process;
 
end project_tb_arch;
